///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: data_source.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::IGLOO> <Die::AGLN250V2> <Package::100 VQFP>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

module data_source( clock, reset, trigger, output_data, tag_control_sig );
input clock, reset;
input trigger;
output reg[19:0] output_data;
output reg[19:0] tag_control_sig;

reg[7:0] tag_data_buf_1;
reg[7:0] tag_data_buf_2;
reg[7:0] tag_data_buf_3;
reg[7:0] tag_data_buf_4;
reg[7:0] tag_data_buf_5;
reg[7:0] tag_data_buf_6;
reg[7:0] tag_data_buf_7;
reg[7:0] tag_data_buf_8;
reg[7:0] tag_data_buf_9;
reg[7:0] tag_data_buf_10;
reg[7:0] tag_data_buf_11;
reg[7:0] tag_data_buf_12;
reg[7:0] tag_data_buf_13;
reg[7:0] tag_data_buf_14;
reg[7:0] tag_data_buf_15;
reg[7:0] tag_data_buf_16;
reg[7:0] tag_data_buf_17;
reg[7:0] tag_data_buf_18;
reg[7:0] tag_data_buf_19;
reg[7:0] tag_data_buf_20;

reg [19:0] tag_order_mem [0:649];

reg[15:0] counter;

always @(posedge clock or negedge reset)
begin
    if (!reset)
    begin
        output_data <= 0;

        tag_data_buf_1 <= 8'd1;
        tag_data_buf_2 <= 8'd2;
        tag_data_buf_3 <= 8'd3;
        tag_data_buf_4 <= 8'd4;
        tag_data_buf_5 <= 8'd5;
        tag_data_buf_6 <= 8'd6;
        tag_data_buf_7 <= 8'd7;
        tag_data_buf_8 <= 8'd8;
        tag_data_buf_9 <= 8'd9;
        tag_data_buf_10 <= 8'd10;
        tag_data_buf_11 <= 8'd11;
        tag_data_buf_12 <= 8'd12;
        tag_data_buf_13 <= 8'd13;
        tag_data_buf_14 <= 8'd14;
        tag_data_buf_15 <= 8'd15;
        tag_data_buf_16 <= 8'd16;
        tag_data_buf_17 <= 8'd17;
        tag_data_buf_18 <= 8'd18;
        tag_data_buf_19 <= 8'd19;
        tag_data_buf_20 <= 8'd20;

        tag_order_mem[0]<=20'd131072;
tag_order_mem[1]<=20'd4098;
tag_order_mem[2]<=20'd16384;
tag_order_mem[3]<=20'd0;
tag_order_mem[4]<=20'd16;
tag_order_mem[5]<=20'd0;
tag_order_mem[6]<=20'd0;
tag_order_mem[7]<=20'd524288;
tag_order_mem[8]<=20'd0;
tag_order_mem[9]<=20'd0;
tag_order_mem[10]<=20'd0;
tag_order_mem[11]<=20'd0;
tag_order_mem[12]<=20'd0;
tag_order_mem[13]<=20'd262240;
tag_order_mem[14]<=20'd512;
tag_order_mem[15]<=20'd33792;
tag_order_mem[16]<=20'd128;
tag_order_mem[17]<=20'd8200;
tag_order_mem[18]<=20'd1;
tag_order_mem[19]<=20'd0;
tag_order_mem[20]<=20'd65536;
tag_order_mem[21]<=20'd0;
tag_order_mem[22]<=20'd0;
tag_order_mem[23]<=20'd4;
tag_order_mem[24]<=20'd2048;
tag_order_mem[25]<=20'd256;
tag_order_mem[26]<=20'd262144;
tag_order_mem[27]<=20'd68;
tag_order_mem[28]<=20'd0;
tag_order_mem[29]<=20'd0;
tag_order_mem[30]<=20'd32;
tag_order_mem[31]<=20'd0;
tag_order_mem[32]<=20'd0;
tag_order_mem[33]<=20'd8192;
tag_order_mem[34]<=20'd0;
tag_order_mem[35]<=20'd0;
tag_order_mem[36]<=20'd0;
tag_order_mem[37]<=20'd256;
tag_order_mem[38]<=20'd0;
tag_order_mem[39]<=20'd0;
tag_order_mem[40]<=20'd0;
tag_order_mem[41]<=20'd2;
tag_order_mem[42]<=20'd0;
tag_order_mem[43]<=20'd1;
tag_order_mem[44]<=20'd16384;
tag_order_mem[45]<=20'd512;
tag_order_mem[46]<=20'd0;
tag_order_mem[47]<=20'd131072;
tag_order_mem[48]<=20'd67584;
tag_order_mem[49]<=20'd557064;
tag_order_mem[50]<=20'd1040;
tag_order_mem[51]<=20'd4224;
tag_order_mem[52]<=20'd0;
tag_order_mem[53]<=20'd65536;
tag_order_mem[54]<=20'd8192;
tag_order_mem[55]<=20'd32;
tag_order_mem[56]<=20'd0;
tag_order_mem[57]<=20'd0;
tag_order_mem[58]<=20'd512;
tag_order_mem[59]<=20'd0;
tag_order_mem[60]<=20'd0;
tag_order_mem[61]<=20'd0;
tag_order_mem[62]<=20'd131072;
tag_order_mem[63]<=20'd0;
tag_order_mem[64]<=20'd32768;
tag_order_mem[65]<=20'd16648;
tag_order_mem[66]<=20'd2;
tag_order_mem[67]<=20'd128;
tag_order_mem[68]<=20'd4097;
tag_order_mem[69]<=20'd64;
tag_order_mem[70]<=20'd0;
tag_order_mem[71]<=20'd4;
tag_order_mem[72]<=20'd786432;
tag_order_mem[73]<=20'd0;
tag_order_mem[74]<=20'd16;
tag_order_mem[75]<=20'd2048;
tag_order_mem[76]<=20'd0;
tag_order_mem[77]<=20'd1024;
tag_order_mem[78]<=20'd32;
tag_order_mem[79]<=20'd0;
tag_order_mem[80]<=20'd0;
tag_order_mem[81]<=20'd1;
tag_order_mem[82]<=20'd0;
tag_order_mem[83]<=20'd0;
tag_order_mem[84]<=20'd4104;
tag_order_mem[85]<=20'd2048;
tag_order_mem[86]<=20'd0;
tag_order_mem[87]<=20'd512;
tag_order_mem[88]<=20'd2;
tag_order_mem[89]<=20'd0;
tag_order_mem[90]<=20'd1024;
tag_order_mem[91]<=20'd0;
tag_order_mem[92]<=20'd32768;
tag_order_mem[93]<=20'd278544;
tag_order_mem[94]<=20'd0;
tag_order_mem[95]<=20'd64;
tag_order_mem[96]<=20'd256;
tag_order_mem[97]<=20'd139264;
tag_order_mem[98]<=20'd524292;
tag_order_mem[99]<=20'd128;
tag_order_mem[100]<=20'd0;
tag_order_mem[101]<=20'd0;
tag_order_mem[102]<=20'd0;
tag_order_mem[103]<=20'd65536;
tag_order_mem[104]<=20'd0;
tag_order_mem[105]<=20'd2;
tag_order_mem[106]<=20'd16384;
tag_order_mem[107]<=20'd0;
tag_order_mem[108]<=20'd0;
tag_order_mem[109]<=20'd270336;
tag_order_mem[110]<=20'd32;
tag_order_mem[111]<=20'd0;
tag_order_mem[112]<=20'd557056;
tag_order_mem[113]<=20'd5248;
tag_order_mem[114]<=20'd16;
tag_order_mem[115]<=20'd0;
tag_order_mem[116]<=20'd4;
tag_order_mem[117]<=20'd0;
tag_order_mem[118]<=20'd65;
tag_order_mem[119]<=20'd0;
tag_order_mem[120]<=20'd131072;
tag_order_mem[121]<=20'd0;
tag_order_mem[122]<=20'd0;
tag_order_mem[123]<=20'd768;
tag_order_mem[124]<=20'd0;
tag_order_mem[125]<=20'd0;
tag_order_mem[126]<=20'd8;
tag_order_mem[127]<=20'd0;
tag_order_mem[128]<=20'd65536;
tag_order_mem[129]<=20'd2048;
tag_order_mem[130]<=20'd0;
tag_order_mem[131]<=20'd262400;
tag_order_mem[132]<=20'd512;
tag_order_mem[133]<=20'd0;
tag_order_mem[134]<=20'd0;
tag_order_mem[135]<=20'd64;
tag_order_mem[136]<=20'd524288;
tag_order_mem[137]<=20'd0;
tag_order_mem[138]<=20'd9217;
tag_order_mem[139]<=20'd32;
tag_order_mem[140]<=20'd0;
tag_order_mem[141]<=20'd16384;
tag_order_mem[142]<=20'd4096;
tag_order_mem[143]<=20'd4;
tag_order_mem[144]<=20'd65544;
tag_order_mem[145]<=20'd0;
tag_order_mem[146]<=20'd0;
tag_order_mem[147]<=20'd32768;
tag_order_mem[148]<=20'd0;
tag_order_mem[149]<=20'd0;
tag_order_mem[150]<=20'd16;
tag_order_mem[151]<=20'd131200;
tag_order_mem[152]<=20'd2048;
tag_order_mem[153]<=20'd2;
tag_order_mem[154]<=20'd0;
tag_order_mem[155]<=20'd0;
tag_order_mem[156]<=20'd0;
tag_order_mem[157]<=20'd8;
tag_order_mem[158]<=20'd131072;
tag_order_mem[159]<=20'd0;
tag_order_mem[160]<=20'd0;
tag_order_mem[161]<=20'd0;
tag_order_mem[162]<=20'd128;
tag_order_mem[163]<=20'd528384;
tag_order_mem[164]<=20'd20;
tag_order_mem[165]<=20'd0;
tag_order_mem[166]<=20'd0;
tag_order_mem[167]<=20'd34;
tag_order_mem[168]<=20'd0;
tag_order_mem[169]<=20'd16384;
tag_order_mem[170]<=20'd2048;
tag_order_mem[171]<=20'd32768;
tag_order_mem[172]<=20'd64;
tag_order_mem[173]<=20'd65537;
tag_order_mem[174]<=20'd262144;
tag_order_mem[175]<=20'd0;
tag_order_mem[176]<=20'd8192;
tag_order_mem[177]<=20'd256;
tag_order_mem[178]<=20'd512;
tag_order_mem[179]<=20'd0;
tag_order_mem[180]<=20'd1024;
tag_order_mem[181]<=20'd0;
tag_order_mem[182]<=20'd2048;
tag_order_mem[183]<=20'd512;
tag_order_mem[184]<=20'd0;
tag_order_mem[185]<=20'd16;
tag_order_mem[186]<=20'd0;
tag_order_mem[187]<=20'd0;
tag_order_mem[188]<=20'd4233;
tag_order_mem[189]<=20'd663620;
tag_order_mem[190]<=20'd2;
tag_order_mem[191]<=20'd0;
tag_order_mem[192]<=20'd0;
tag_order_mem[193]<=20'd0;
tag_order_mem[194]<=20'd0;
tag_order_mem[195]<=20'd0;
tag_order_mem[196]<=20'd256;
tag_order_mem[197]<=20'd0;
tag_order_mem[198]<=20'd32768;
tag_order_mem[199]<=20'd16416;
tag_order_mem[200]<=20'd65536;
tag_order_mem[201]<=20'd0;
tag_order_mem[202]<=20'd0;
tag_order_mem[203]<=20'd1024;
tag_order_mem[204]<=20'd0;
tag_order_mem[205]<=20'd0;
tag_order_mem[206]<=20'd0;
tag_order_mem[207]<=20'd262144;
tag_order_mem[208]<=20'd0;
tag_order_mem[209]<=20'd49168;
tag_order_mem[210]<=20'd0;
tag_order_mem[211]<=20'd8194;
tag_order_mem[212]<=20'd0;
tag_order_mem[213]<=20'd128;
tag_order_mem[214]<=20'd8;
tag_order_mem[215]<=20'd256;
tag_order_mem[216]<=20'd0;
tag_order_mem[217]<=20'd32;
tag_order_mem[218]<=20'd2048;
tag_order_mem[219]<=20'd0;
tag_order_mem[220]<=20'd0;
tag_order_mem[221]<=20'd524801;
tag_order_mem[222]<=20'd65536;
tag_order_mem[223]<=20'd262144;
tag_order_mem[224]<=20'd1024;
tag_order_mem[225]<=20'd4096;
tag_order_mem[226]<=20'd0;
tag_order_mem[227]<=20'd0;
tag_order_mem[228]<=20'd0;
tag_order_mem[229]<=20'd0;
tag_order_mem[230]<=20'd0;
tag_order_mem[231]<=20'd131076;
tag_order_mem[232]<=20'd0;
tag_order_mem[233]<=20'd64;
tag_order_mem[234]<=20'd256;
tag_order_mem[235]<=20'd262144;
tag_order_mem[236]<=20'd65536;
tag_order_mem[237]<=20'd0;
tag_order_mem[238]<=20'd0;
tag_order_mem[239]<=20'd0;
tag_order_mem[240]<=20'd68;
tag_order_mem[241]<=20'd640;
tag_order_mem[242]<=20'd0;
tag_order_mem[243]<=20'd1024;
tag_order_mem[244]<=20'd2;
tag_order_mem[245]<=20'd0;
tag_order_mem[246]<=20'd0;
tag_order_mem[247]<=20'd131072;
tag_order_mem[248]<=20'd0;
tag_order_mem[249]<=20'd4104;
tag_order_mem[250]<=20'd2065;
tag_order_mem[251]<=20'd0;
tag_order_mem[252]<=20'd0;
tag_order_mem[253]<=20'd8224;
tag_order_mem[254]<=20'd524288;
tag_order_mem[255]<=20'd0;
tag_order_mem[256]<=20'd16384;
tag_order_mem[257]<=20'd32768;
tag_order_mem[258]<=20'd0;
tag_order_mem[259]<=20'd0;
tag_order_mem[260]<=20'd0;
tag_order_mem[261]<=20'd1024;
tag_order_mem[262]<=20'd512;
tag_order_mem[263]<=20'd8;
tag_order_mem[264]<=20'd0;
tag_order_mem[265]<=20'd32784;
tag_order_mem[266]<=20'd262;
tag_order_mem[267]<=20'd133120;
tag_order_mem[268]<=20'd1;
tag_order_mem[269]<=20'd0;
tag_order_mem[270]<=20'd65536;
tag_order_mem[271]<=20'd0;
tag_order_mem[272]<=20'd0;
tag_order_mem[273]<=20'd0;
tag_order_mem[274]<=20'd16384;
tag_order_mem[275]<=20'd0;
tag_order_mem[276]<=20'd8192;
tag_order_mem[277]<=20'd4096;
tag_order_mem[278]<=20'd0;
tag_order_mem[279]<=20'd524480;
tag_order_mem[280]<=20'd0;
tag_order_mem[281]<=20'd262176;
tag_order_mem[282]<=20'd0;
tag_order_mem[283]<=20'd0;
tag_order_mem[284]<=20'd0;
tag_order_mem[285]<=20'd0;
tag_order_mem[286]<=20'd0;
tag_order_mem[287]<=20'd131080;
tag_order_mem[288]<=20'd0;
tag_order_mem[289]<=20'd8192;
tag_order_mem[290]<=20'd0;
tag_order_mem[291]<=20'd0;
tag_order_mem[292]<=20'd544832;
tag_order_mem[293]<=20'd0;
tag_order_mem[294]<=20'd1024;
tag_order_mem[295]<=20'd32768;
tag_order_mem[296]<=20'd2;
tag_order_mem[297]<=20'd0;
tag_order_mem[298]<=20'd256;
tag_order_mem[299]<=20'd0;
tag_order_mem[300]<=20'd2048;
tag_order_mem[301]<=20'd0;
tag_order_mem[302]<=20'd0;
tag_order_mem[303]<=20'd327712;
tag_order_mem[304]<=20'd0;
tag_order_mem[305]<=20'd132;
tag_order_mem[306]<=20'd0;
tag_order_mem[307]<=20'd0;
tag_order_mem[308]<=20'd513;
tag_order_mem[309]<=20'd0;
tag_order_mem[310]<=20'd16;
tag_order_mem[311]<=20'd0;
tag_order_mem[312]<=20'd0;
tag_order_mem[313]<=20'd16384;
tag_order_mem[314]<=20'd0;
tag_order_mem[315]<=20'd264;
tag_order_mem[316]<=20'd0;
tag_order_mem[317]<=20'd32768;
tag_order_mem[318]<=20'd16;
tag_order_mem[319]<=20'd4096;
tag_order_mem[320]<=20'd0;
tag_order_mem[321]<=20'd0;
tag_order_mem[322]<=20'd32;
tag_order_mem[323]<=20'd1028;
tag_order_mem[324]<=20'd0;
tag_order_mem[325]<=20'd128;
tag_order_mem[326]<=20'd2;
tag_order_mem[327]<=20'd524288;
tag_order_mem[328]<=20'd0;
tag_order_mem[329]<=20'd0;
tag_order_mem[330]<=20'd131072;
tag_order_mem[331]<=20'd0;
tag_order_mem[332]<=20'd73728;
tag_order_mem[333]<=20'd0;
tag_order_mem[334]<=20'd1;
tag_order_mem[335]<=20'd264704;
tag_order_mem[336]<=20'd0;
tag_order_mem[337]<=20'd64;
tag_order_mem[338]<=20'd512;
tag_order_mem[339]<=20'd128;
tag_order_mem[340]<=20'd0;
tag_order_mem[341]<=20'd16384;
tag_order_mem[342]<=20'd0;
tag_order_mem[343]<=20'd131072;
tag_order_mem[344]<=20'd524544;
tag_order_mem[345]<=20'd4096;
tag_order_mem[346]<=20'd32768;
tag_order_mem[347]<=20'd1024;
tag_order_mem[348]<=20'd65600;
tag_order_mem[349]<=20'd0;
tag_order_mem[350]<=20'd0;
tag_order_mem[351]<=20'd0;
tag_order_mem[352]<=20'd1;
tag_order_mem[353]<=20'd0;
tag_order_mem[354]<=20'd0;
tag_order_mem[355]<=20'd32;
tag_order_mem[356]<=20'd0;
tag_order_mem[357]<=20'd262146;
tag_order_mem[358]<=20'd0;
tag_order_mem[359]<=20'd0;
tag_order_mem[360]<=20'd8212;
tag_order_mem[361]<=20'd2056;
tag_order_mem[362]<=20'd0;
tag_order_mem[363]<=20'd0;
tag_order_mem[364]<=20'd0;
tag_order_mem[365]<=20'd0;
tag_order_mem[366]<=20'd0;
tag_order_mem[367]<=20'd0;
tag_order_mem[368]<=20'd4;
tag_order_mem[369]<=20'd1024;
tag_order_mem[370]<=20'd69632;
tag_order_mem[371]<=20'd2;
tag_order_mem[372]<=20'd0;
tag_order_mem[373]<=20'd0;
tag_order_mem[374]<=20'd0;
tag_order_mem[375]<=20'd8192;
tag_order_mem[376]<=20'd0;
tag_order_mem[377]<=20'd0;
tag_order_mem[378]<=20'd0;
tag_order_mem[379]<=20'd0;
tag_order_mem[380]<=20'd2048;
tag_order_mem[381]<=20'd0;
tag_order_mem[382]<=20'd32840;
tag_order_mem[383]<=20'd131072;
tag_order_mem[384]<=20'd16384;
tag_order_mem[385]<=20'd524416;
tag_order_mem[386]<=20'd256;
tag_order_mem[387]<=20'd262689;
tag_order_mem[388]<=20'd16;
tag_order_mem[389]<=20'd0;
tag_order_mem[390]<=20'd131072;
tag_order_mem[391]<=20'd0;
tag_order_mem[392]<=20'd128;
tag_order_mem[393]<=20'd514;
tag_order_mem[394]<=20'd0;
tag_order_mem[395]<=20'd73728;
tag_order_mem[396]<=20'd0;
tag_order_mem[397]<=20'd1024;
tag_order_mem[398]<=20'd524288;
tag_order_mem[399]<=20'd2112;
tag_order_mem[400]<=20'd32768;
tag_order_mem[401]<=20'd288;
tag_order_mem[402]<=20'd0;
tag_order_mem[403]<=20'd0;
tag_order_mem[404]<=20'd0;
tag_order_mem[405]<=20'd0;
tag_order_mem[406]<=20'd0;
tag_order_mem[407]<=20'd16384;
tag_order_mem[408]<=20'd0;
tag_order_mem[409]<=20'd24;
tag_order_mem[410]<=20'd262144;
tag_order_mem[411]<=20'd0;
tag_order_mem[412]<=20'd4;
tag_order_mem[413]<=20'd0;
tag_order_mem[414]<=20'd4096;
tag_order_mem[415]<=20'd1;
tag_order_mem[416]<=20'd512;
tag_order_mem[417]<=20'd0;
tag_order_mem[418]<=20'd2048;
tag_order_mem[419]<=20'd4096;
tag_order_mem[420]<=20'd0;
tag_order_mem[421]<=20'd147456;
tag_order_mem[422]<=20'd0;
tag_order_mem[423]<=20'd4;
tag_order_mem[424]<=20'd0;
tag_order_mem[425]<=20'd0;
tag_order_mem[426]<=20'd0;
tag_order_mem[427]<=20'd0;
tag_order_mem[428]<=20'd0;
tag_order_mem[429]<=20'd0;
tag_order_mem[430]<=20'd128;
tag_order_mem[431]<=20'd524322;
tag_order_mem[432]<=20'd0;
tag_order_mem[433]<=20'd0;
tag_order_mem[434]<=20'd270336;
tag_order_mem[435]<=20'd32769;
tag_order_mem[436]<=20'd0;
tag_order_mem[437]<=20'd328;
tag_order_mem[438]<=20'd66560;
tag_order_mem[439]<=20'd16;
tag_order_mem[440]<=20'd0;
tag_order_mem[441]<=20'd0;
tag_order_mem[442]<=20'd65792;
tag_order_mem[443]<=20'd2048;
tag_order_mem[444]<=20'd0;
tag_order_mem[445]<=20'd4096;
tag_order_mem[446]<=20'd4;
tag_order_mem[447]<=20'd8;
tag_order_mem[448]<=20'd139264;
tag_order_mem[449]<=20'd0;
tag_order_mem[450]<=20'd512;
tag_order_mem[451]<=20'd64;
tag_order_mem[452]<=20'd0;
tag_order_mem[453]<=20'd0;
tag_order_mem[454]<=20'd0;
tag_order_mem[455]<=20'd1;
tag_order_mem[456]<=20'd0;
tag_order_mem[457]<=20'd262144;
tag_order_mem[458]<=20'd1024;
tag_order_mem[459]<=20'd16;
tag_order_mem[460]<=20'd0;
tag_order_mem[461]<=20'd32;
tag_order_mem[462]<=20'd0;
tag_order_mem[463]<=20'd0;
tag_order_mem[464]<=20'd16384;
tag_order_mem[465]<=20'd32768;
tag_order_mem[466]<=20'd2;
tag_order_mem[467]<=20'd524416;
tag_order_mem[468]<=20'd0;
tag_order_mem[469]<=20'd0;
tag_order_mem[470]<=20'd0;
tag_order_mem[471]<=20'd24576;
tag_order_mem[472]<=20'd0;
tag_order_mem[473]<=20'd16;
tag_order_mem[474]<=20'd4096;
tag_order_mem[475]<=20'd128;
tag_order_mem[476]<=20'd65536;
tag_order_mem[477]<=20'd8;
tag_order_mem[478]<=20'd0;
tag_order_mem[479]<=20'd0;
tag_order_mem[480]<=20'd0;
tag_order_mem[481]<=20'd0;
tag_order_mem[482]<=20'd96;
tag_order_mem[483]<=20'd0;
tag_order_mem[484]<=20'd132098;
tag_order_mem[485]<=20'd32768;
tag_order_mem[486]<=20'd2048;
tag_order_mem[487]<=20'd524288;
tag_order_mem[488]<=20'd262144;
tag_order_mem[489]<=20'd512;
tag_order_mem[490]<=20'd256;
tag_order_mem[491]<=20'd0;
tag_order_mem[492]<=20'd4;
tag_order_mem[493]<=20'd1;
tag_order_mem[494]<=20'd1024;
tag_order_mem[495]<=20'd32834;
tag_order_mem[496]<=20'd65536;
tag_order_mem[497]<=20'd0;
tag_order_mem[498]<=20'd0;
tag_order_mem[499]<=20'd4;
tag_order_mem[500]<=20'd4096;
tag_order_mem[501]<=20'd0;
tag_order_mem[502]<=20'd0;
tag_order_mem[503]<=20'd655360;
tag_order_mem[504]<=20'd0;
tag_order_mem[505]<=20'd16384;
tag_order_mem[506]<=20'd8;
tag_order_mem[507]<=20'd262656;
tag_order_mem[508]<=20'd32;
tag_order_mem[509]<=20'd0;
tag_order_mem[510]<=20'd0;
tag_order_mem[511]<=20'd0;
tag_order_mem[512]<=20'd0;
tag_order_mem[513]<=20'd1;
tag_order_mem[514]<=20'd384;
tag_order_mem[515]<=20'd0;
tag_order_mem[516]<=20'd0;
tag_order_mem[517]<=20'd8208;
tag_order_mem[518]<=20'd0;
tag_order_mem[519]<=20'd2048;
tag_order_mem[520]<=20'd1;
tag_order_mem[521]<=20'd65536;
tag_order_mem[522]<=20'd2048;
tag_order_mem[523]<=20'd0;
tag_order_mem[524]<=20'd1296;
tag_order_mem[525]<=20'd0;
tag_order_mem[526]<=20'd147456;
tag_order_mem[527]<=20'd0;
tag_order_mem[528]<=20'd4;
tag_order_mem[529]<=20'd0;
tag_order_mem[530]<=20'd0;
tag_order_mem[531]<=20'd64;
tag_order_mem[532]<=20'd0;
tag_order_mem[533]<=20'd0;
tag_order_mem[534]<=20'd0;
tag_order_mem[535]<=20'd32768;
tag_order_mem[536]<=20'd32;
tag_order_mem[537]<=20'd524424;
tag_order_mem[538]<=20'd2;
tag_order_mem[539]<=20'd4096;
tag_order_mem[540]<=20'd0;
tag_order_mem[541]<=20'd0;
tag_order_mem[542]<=20'd262144;
tag_order_mem[543]<=20'd8704;
tag_order_mem[544]<=20'd0;
tag_order_mem[545]<=20'd0;
tag_order_mem[546]<=20'd0;
tag_order_mem[547]<=20'd512;
tag_order_mem[548]<=20'd256;
tag_order_mem[549]<=20'd393216;
tag_order_mem[550]<=20'd0;
tag_order_mem[551]<=20'd12;
tag_order_mem[552]<=20'd65536;
tag_order_mem[553]<=20'd0;
tag_order_mem[554]<=20'd0;
tag_order_mem[555]<=20'd2;
tag_order_mem[556]<=20'd32;
tag_order_mem[557]<=20'd0;
tag_order_mem[558]<=20'd8193;
tag_order_mem[559]<=20'd128;
tag_order_mem[560]<=20'd32768;
tag_order_mem[561]<=20'd2048;
tag_order_mem[562]<=20'd0;
tag_order_mem[563]<=20'd0;
tag_order_mem[564]<=20'd0;
tag_order_mem[565]<=20'd524304;
tag_order_mem[566]<=20'd0;
tag_order_mem[567]<=20'd64;
tag_order_mem[568]<=20'd0;
tag_order_mem[569]<=20'd0;
tag_order_mem[570]<=20'd1024;
tag_order_mem[571]<=20'd20480;
tag_order_mem[572]<=20'd0;
tag_order_mem[573]<=20'd32768;
tag_order_mem[574]<=20'd32;
tag_order_mem[575]<=20'd1;
tag_order_mem[576]<=20'd16450;
tag_order_mem[577]<=20'd0;
tag_order_mem[578]<=20'd0;
tag_order_mem[579]<=20'd1024;
tag_order_mem[580]<=20'd8;
tag_order_mem[581]<=20'd512;
tag_order_mem[582]<=20'd139268;
tag_order_mem[583]<=20'd16;
tag_order_mem[584]<=20'd0;
tag_order_mem[585]<=20'd524288;
tag_order_mem[586]<=20'd0;
tag_order_mem[587]<=20'd262144;
tag_order_mem[588]<=20'd128;
tag_order_mem[589]<=20'd0;
tag_order_mem[590]<=20'd4096;
tag_order_mem[591]<=20'd0;
tag_order_mem[592]<=20'd256;
tag_order_mem[593]<=20'd0;
tag_order_mem[594]<=20'd0;
tag_order_mem[595]<=20'd2048;
tag_order_mem[596]<=20'd65536;
tag_order_mem[597]<=20'd0;
tag_order_mem[598]<=20'd0;
tag_order_mem[599]<=20'd24;
tag_order_mem[600]<=20'd4;
tag_order_mem[601]<=20'd0;
tag_order_mem[602]<=20'd2;
tag_order_mem[603]<=20'd0;
tag_order_mem[604]<=20'd0;
tag_order_mem[605]<=20'd524288;
tag_order_mem[606]<=20'd0;
tag_order_mem[607]<=20'd0;
tag_order_mem[608]<=20'd256;
tag_order_mem[609]<=20'd8192;
tag_order_mem[610]<=20'd69696;
tag_order_mem[611]<=20'd49152;
tag_order_mem[612]<=20'd0;
tag_order_mem[613]<=20'd0;
tag_order_mem[614]<=20'd0;
tag_order_mem[615]<=20'd32;
tag_order_mem[616]<=20'd1024;
tag_order_mem[617]<=20'd0;
tag_order_mem[618]<=20'd0;
tag_order_mem[619]<=20'd0;
tag_order_mem[620]<=20'd262656;
tag_order_mem[621]<=20'd1;
tag_order_mem[622]<=20'd133248;
tag_order_mem[623]<=20'd0;
tag_order_mem[624]<=20'd0;
tag_order_mem[625]<=20'd131072;
tag_order_mem[626]<=20'd16;
tag_order_mem[627]<=20'd262144;
tag_order_mem[628]<=20'd8;
tag_order_mem[629]<=20'd512;
tag_order_mem[630]<=20'd16384;
tag_order_mem[631]<=20'd1028;
tag_order_mem[632]<=20'd0;
tag_order_mem[633]<=20'd0;
tag_order_mem[634]<=20'd8192;
tag_order_mem[635]<=20'd4224;
tag_order_mem[636]<=20'd524288;
tag_order_mem[637]<=20'd64;
tag_order_mem[638]<=20'd0;
tag_order_mem[639]<=20'd32768;
tag_order_mem[640]<=20'd0;
tag_order_mem[641]<=20'd0;
tag_order_mem[642]<=20'd1;
tag_order_mem[643]<=20'd2080;
tag_order_mem[644]<=20'd256;
tag_order_mem[645]<=20'd65536;
tag_order_mem[646]<=20'd2;
tag_order_mem[647]<=20'd0;
tag_order_mem[648]<=20'd0;
tag_order_mem[649]<=20'd0;

        counter <= 0;
    end
    else if (trigger)
    begin
        if (counter==16'd0)
        begin
            counter <= counter+1;
            tag_data_buf_1 <= {tag_data_buf_1[6:0],tag_data_buf_1[7]};
            tag_data_buf_2 <= {tag_data_buf_2[6:0],tag_data_buf_2[7]};
            tag_data_buf_3 <= {tag_data_buf_3[6:0],tag_data_buf_3[7]};
            tag_data_buf_4 <= {tag_data_buf_4[6:0],tag_data_buf_4[7]};
            tag_data_buf_5 <= {tag_data_buf_5[6:0],tag_data_buf_5[7]};
            tag_data_buf_6 <= {tag_data_buf_6[6:0],tag_data_buf_6[7]};
            tag_data_buf_7 <= {tag_data_buf_7[6:0],tag_data_buf_7[7]};
            tag_data_buf_8 <= {tag_data_buf_8[6:0],tag_data_buf_8[7]};
            tag_data_buf_9 <= {tag_data_buf_9[6:0],tag_data_buf_9[7]};
            tag_data_buf_10 <= {tag_data_buf_10[6:0],tag_data_buf_10[7]};
            tag_data_buf_11 <= {tag_data_buf_11[6:0],tag_data_buf_11[7]};
            tag_data_buf_12 <= {tag_data_buf_12[6:0],tag_data_buf_12[7]};
            tag_data_buf_13 <= {tag_data_buf_13[6:0],tag_data_buf_13[7]};
            tag_data_buf_14 <= {tag_data_buf_14[6:0],tag_data_buf_14[7]};
            tag_data_buf_15 <= {tag_data_buf_15[6:0],tag_data_buf_15[7]};
            tag_data_buf_16 <= {tag_data_buf_16[6:0],tag_data_buf_16[7]};
            tag_data_buf_17 <= {tag_data_buf_17[6:0],tag_data_buf_17[7]};
            tag_data_buf_18 <= {tag_data_buf_18[6:0],tag_data_buf_18[7]};
            tag_data_buf_19 <= {tag_data_buf_19[6:0],tag_data_buf_19[7]};
            tag_data_buf_20 <= {tag_data_buf_20[6:0],tag_data_buf_20[7]};

            output_data[0] <= tag_data_buf_1[7];
            output_data[1] <= tag_data_buf_2[7];
            output_data[2] <= tag_data_buf_3[7];
            output_data[3] <= tag_data_buf_4[7];
            output_data[4] <= tag_data_buf_5[7];
            output_data[5] <= tag_data_buf_6[7];
            output_data[6] <= tag_data_buf_7[7];
            output_data[7] <= tag_data_buf_8[7];
            output_data[8] <= tag_data_buf_9[7];
            output_data[9] <= tag_data_buf_10[7];
            output_data[10] <= tag_data_buf_11[7];
            output_data[11] <= tag_data_buf_12[7];
            output_data[12] <= tag_data_buf_13[7];
            output_data[13] <= tag_data_buf_14[7];
            output_data[14] <= tag_data_buf_15[7];
            output_data[15] <= tag_data_buf_16[7];
            output_data[16] <= tag_data_buf_17[7];
            output_data[17] <= tag_data_buf_18[7];
            output_data[18] <= tag_data_buf_19[7];
            output_data[19] <= tag_data_buf_20[7];
        end
        else
        begin
            counter <= counter + 1;
            if (counter==16'd799)
                counter <= 0;
        end
    end
    else
    begin
        output_data <= 0;

        tag_data_buf_1 <= 8'd1;
        tag_data_buf_2 <= 8'd2;
        tag_data_buf_3 <= 8'd3;
        tag_data_buf_4 <= 8'd4;
        tag_data_buf_5 <= 8'd5;
        tag_data_buf_6 <= 8'd6;
        tag_data_buf_7 <= 8'd7;
        tag_data_buf_8 <= 8'd8;
        tag_data_buf_9 <= 8'd9;
        tag_data_buf_10 <= 8'd10;
        tag_data_buf_11 <= 8'd11;
        tag_data_buf_12 <= 8'd12;
        tag_data_buf_13 <= 8'd13;
        tag_data_buf_14 <= 8'd14;
        tag_data_buf_15 <= 8'd15;
        tag_data_buf_16 <= 8'd16;
        tag_data_buf_17 <= 8'd17;
        tag_data_buf_18 <= 8'd18;
        tag_data_buf_19 <= 8'd19;
        tag_data_buf_20 <= 8'd20;

        tag_control_sig <= tag_order_mem[data_index];

        counter <= 0;
    end
end

reg[16:0] data_index;
reg[7:0] trigger_counter;

always @(posedge trigger or negedge reset)
begin
    if (!reset)
    begin
        data_index <= 1;
        trigger_counter <= 0;
    end
    else
    begin
        //trigger_counter <= trigger_counter+1;
        //if(trigger_counter==8'd9)
        begin
            //trigger_counter <= 0;
            if(data_index<=16'd648)
                data_index <= data_index + 1;
            else
                data_index <= 16'd0;
        end
    end
end

endmodule

