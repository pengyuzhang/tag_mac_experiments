`timescale 1 ns/100 ps
// Version: v11.8 11.8.0.26
// File used only for Simulation


module PLLBA(
       CLKA,
       EXTFB,
       POWERDOWN,
       GLA,
       LOCK,
       GLB,
       YB,
       GLC,
       YC,
       OADIV0,
       OADIV1,
       OADIV2,
       OADIV3,
       OADIV4,
       OAMUX0,
       OAMUX1,
       OAMUX2,
       DLYGLA0,
       DLYGLA1,
       DLYGLA2,
       DLYGLA3,
       DLYGLA4,
       OBDIV0,
       OBDIV1,
       OBDIV2,
       OBDIV3,
       OBDIV4,
       OBMUX0,
       OBMUX1,
       OBMUX2,
       DLYYB0,
       DLYYB1,
       DLYYB2,
       DLYYB3,
       DLYYB4,
       DLYGLB0,
       DLYGLB1,
       DLYGLB2,
       DLYGLB3,
       DLYGLB4,
       OCDIV0,
       OCDIV1,
       OCDIV2,
       OCDIV3,
       OCDIV4,
       OCMUX0,
       OCMUX1,
       OCMUX2,
       DLYYC0,
       DLYYC1,
       DLYYC2,
       DLYYC3,
       DLYYC4,
       DLYGLC0,
       DLYGLC1,
       DLYGLC2,
       DLYGLC3,
       DLYGLC4,
       FINDIV0,
       FINDIV1,
       FINDIV2,
       FINDIV3,
       FINDIV4,
       FINDIV5,
       FINDIV6,
       FBDIV0,
       FBDIV1,
       FBDIV2,
       FBDIV3,
       FBDIV4,
       FBDIV5,
       FBDIV6,
       FBDLY0,
       FBDLY1,
       FBDLY2,
       FBDLY3,
       FBDLY4,
       FBSEL0,
       FBSEL1,
       XDLYSEL,
       VCOSEL0,
       VCOSEL1,
       VCOSEL2
    );
input  CLKA;
input  EXTFB;
input  POWERDOWN;
output GLA;
output LOCK;
output GLB;
output YB;
output GLC;
output YC;
input  OADIV0;
input  OADIV1;
input  OADIV2;
input  OADIV3;
input  OADIV4;
input  OAMUX0;
input  OAMUX1;
input  OAMUX2;
input  DLYGLA0;
input  DLYGLA1;
input  DLYGLA2;
input  DLYGLA3;
input  DLYGLA4;
input  OBDIV0;
input  OBDIV1;
input  OBDIV2;
input  OBDIV3;
input  OBDIV4;
input  OBMUX0;
input  OBMUX1;
input  OBMUX2;
input  DLYYB0;
input  DLYYB1;
input  DLYYB2;
input  DLYYB3;
input  DLYYB4;
input  DLYGLB0;
input  DLYGLB1;
input  DLYGLB2;
input  DLYGLB3;
input  DLYGLB4;
input  OCDIV0;
input  OCDIV1;
input  OCDIV2;
input  OCDIV3;
input  OCDIV4;
input  OCMUX0;
input  OCMUX1;
input  OCMUX2;
input  DLYYC0;
input  DLYYC1;
input  DLYYC2;
input  DLYYC3;
input  DLYYC4;
input  DLYGLC0;
input  DLYGLC1;
input  DLYGLC2;
input  DLYGLC3;
input  DLYGLC4;
input  FINDIV0;
input  FINDIV1;
input  FINDIV2;
input  FINDIV3;
input  FINDIV4;
input  FINDIV5;
input  FINDIV6;
input  FBDIV0;
input  FBDIV1;
input  FBDIV2;
input  FBDIV3;
input  FBDIV4;
input  FBDIV5;
input  FBDIV6;
input  FBDLY0;
input  FBDLY1;
input  FBDLY2;
input  FBDLY3;
input  FBDLY4;
input  FBSEL0;
input  FBSEL1;
input  XDLYSEL;
input  VCOSEL0;
input  VCOSEL1;
input  VCOSEL2;

    wire GND, SDOUT, FB, EXTFBDLY, GLADLY, LOCKDLY, GLBDLY, YBDLY, 
        GLCDLY, YCDLY, VCODLY;
    wire GND_power_net1;
    assign GND = GND_power_net1;
    
    PLL_SDF #( .VCOFREQUENCY(100.000000) )  pll_sdf_0 (.CLKA(CLKA), 
        .EXTFB(EXTFBDLY), .POWERDOWN(POWERDOWN), .GLAOUT(GLADLY), 
        .LOCKOUT(LOCKDLY), .GLBOUT(GLBDLY), .YBOUT(YBDLY), .GLCOUT(
        GLCDLY), .YCOUT(YCDLY), .OADIV0(OADIV0), .OADIV1(OADIV1), 
        .OADIV2(OADIV2), .OADIV3(OADIV3), .OADIV4(OADIV4), .OAMUX0(
        OAMUX0), .OAMUX1(OAMUX1), .OAMUX2(OAMUX2), .DLYGLA0(DLYGLA0), 
        .DLYGLA1(DLYGLA1), .DLYGLA2(DLYGLA2), .DLYGLA3(DLYGLA3), 
        .DLYGLA4(DLYGLA4), .OBDIV0(OBDIV0), .OBDIV1(OBDIV1), .OBDIV2(
        OBDIV2), .OBDIV3(OBDIV3), .OBDIV4(OBDIV4), .OBMUX0(OBMUX0), 
        .OBMUX1(OBMUX1), .OBMUX2(OBMUX2), .DLYYB0(DLYYB0), .DLYYB1(
        DLYYB1), .DLYYB2(DLYYB2), .DLYYB3(DLYYB3), .DLYYB4(DLYYB4), 
        .DLYGLB0(DLYGLB0), .DLYGLB1(DLYGLB1), .DLYGLB2(DLYGLB2), 
        .DLYGLB3(DLYGLB3), .DLYGLB4(DLYGLB4), .OCDIV0(OCDIV0), .OCDIV1(
        OCDIV1), .OCDIV2(OCDIV2), .OCDIV3(OCDIV3), .OCDIV4(OCDIV4), 
        .OCMUX0(OCMUX0), .OCMUX1(OCMUX1), .OCMUX2(OCMUX2), .DLYYC0(
        DLYYC0), .DLYYC1(DLYYC1), .DLYYC2(DLYYC2), .DLYYC3(DLYYC3), 
        .DLYYC4(DLYYC4), .DLYGLC0(DLYGLC0), .DLYGLC1(DLYGLC1), 
        .DLYGLC2(DLYGLC2), .DLYGLC3(DLYGLC3), .DLYGLC4(DLYGLC4), 
        .FINDIV0(FINDIV0), .FINDIV1(FINDIV1), .FINDIV2(FINDIV2), 
        .FINDIV3(FINDIV3), .FINDIV4(FINDIV4), .FINDIV5(FINDIV5), 
        .FINDIV6(FINDIV6), .FBDIV0(FBDIV0), .FBDIV1(FBDIV1), .FBDIV2(
        FBDIV2), .FBDIV3(FBDIV3), .FBDIV4(FBDIV4), .FBDIV5(FBDIV5), 
        .FBDIV6(FBDIV6), .FBDLY0(FBDLY0), .FBDLY1(FBDLY1), .FBDLY2(
        FBDLY2), .FBDLY3(FBDLY3), .FBDLY4(FBDLY4), .FBSEL0(FBSEL0), 
        .FBSEL1(FBSEL1), .XDLYSEL(XDLYSEL), .VCOSEL0(VCOSEL0), 
        .VCOSEL1(VCOSEL1), .VCOSEL2(VCOSEL2), .INTFB(FB), .VCOOUT(
        VCODLY));
    PLL_DLY_SDF #( .VCOFREQUENCY(100.000000) )  pll_dly_sdf_0 (.GLA(
        GLA), .LOCK(LOCK), .GLB(GLB), .YB(YB), .GLC(GLC), .YC(YC), 
        .GLAIN(GLADLY), .LOCKIN(LOCKDLY), .GLBIN(GLBDLY), .YBIN(YBDLY), 
        .GLCIN(GLCDLY), .YCIN(YCDLY), .EXTFBOUT(EXTFBDLY), .EXTFBIN(
        EXTFB), .VCOIN(VCODLY), .PLLOUT(FB));
    GND GND_power_inst1 (.Y(GND_power_net1));
    
endmodule


module top(
       clock,
       mac_control_signal,
       reset,
       trigger_signal,
       output_signal,
       signal_into_switch
    );
input  clock;
input  mac_control_signal;
input  reset;
input  trigger_signal;
output [19:0] output_signal;
output signal_into_switch;

    wire AND2_0_Y, main_clock_0_clock_out, 
        \data_source_0_output_data_0[0] , 
        \data_source_0_output_data_0[1] , 
        \data_source_0_output_data_0[2] , 
        \data_source_0_output_data_0[3] , 
        \data_source_0_output_data_0[4] , 
        \data_source_0_output_data_0[5] , 
        \data_source_0_output_data_0[6] , 
        \data_source_0_output_data_0[7] , 
        \data_source_0_output_data_0[9] , 
        \data_source_0_output_data_0[10] , 
        \data_source_0_output_data_0[11] , 
        \data_source_0_output_data_0[12] , 
        \data_source_0_output_data_0[13] , 
        \data_source_0_output_data_0[14] , 
        \data_source_0_output_data_0[15] , 
        \data_source_0_output_data_0[16] , 
        \data_source_0_output_data_0[17] , 
        \data_source_0_output_data_0[18] , 
        \data_source_0_output_data_0[19] , modulator_0_output_signal, 
        \data_source_0_tag_control_sig[0] , 
        \data_source_0_tag_control_sig[1] , 
        \data_source_0_tag_control_sig[2] , 
        \data_source_0_tag_control_sig[3] , 
        \data_source_0_tag_control_sig[4] , 
        \data_source_0_tag_control_sig[5] , 
        \data_source_0_tag_control_sig[6] , 
        \data_source_0_tag_control_sig[7] , 
        \data_source_0_tag_control_sig[8] , 
        \data_source_0_tag_control_sig[9] , 
        \data_source_0_tag_control_sig[10] , 
        \data_source_0_tag_control_sig[11] , 
        \data_source_0_tag_control_sig[12] , 
        \data_source_0_tag_control_sig[13] , 
        \data_source_0_tag_control_sig[14] , 
        \data_source_0_tag_control_sig[15] , 
        \data_source_0_tag_control_sig[16] , 
        \data_source_0_tag_control_sig[17] , 
        \data_source_0_tag_control_sig[18] , 
        \data_source_0_tag_control_sig[19] , GLA, clock_c, 
        mac_control_signal_c, reset_c, trigger_signal_c, 
        \output_signal_c[0] , \output_signal_c[1] , 
        \output_signal_c[2] , \output_signal_c[3] , 
        \output_signal_c[4] , \output_signal_c[5] , 
        \output_signal_c[6] , \output_signal_c[7] , 
        \output_signal_c[8] , \output_signal_c[9] , 
        \output_signal_c[10] , \output_signal_c[11] , 
        \output_signal_c[12] , \output_signal_c[13] , 
        \output_signal_c[14] , \output_signal_c[15] , 
        \output_signal_c[16] , \output_signal_c[17] , 
        \output_signal_c[18] , \output_signal_c[19] , 
        \modulator_0/output_signal_i , 
        \modulator_0/clock_counter[14]_net_1 , 
        \modulator_0/output_signal_1_sqmuxa_0 , 
        \modulator_0/un5lto15_5 , \modulator_0/un5lto15_6 , 
        \modulator_0/un6lto15_1 , 
        \modulator_0/clock_counter[13]_net_1 , 
        \modulator_0/clock_counter[15]_net_1 , 
        \modulator_0/un5lto15_2 , \modulator_0/un5lto15_1 , 
        \modulator_0/un5lto15_3 , \modulator_0/un5lto5 , 
        \modulator_0/un5lto6 , \modulator_0/un6lto8 , 
        \modulator_0/un6lto9 , \modulator_0/un6lto10 , 
        \modulator_0/un6lto12 , \modulator_0/un6lto11 , 
        \modulator_0/un6lto6_0 , \modulator_0/clock_counter[5]_net_1 , 
        \modulator_0/counter19_1 , \modulator_0/counter[4]_net_1 , 
        \modulator_0/counter[0]_net_1 , \modulator_0/counter19_0 , 
        \modulator_0/counter[5]_net_1 , \modulator_0/counter[1]_net_1 , 
        \modulator_0/un6lt4_2 , \modulator_0/clock_counter[0]_net_1 , 
        \modulator_0/clock_counter[1]_net_1 , 
        \modulator_0/clock_counter[4]_net_1 , 
        \modulator_0/counter23_2 , \modulator_0/counter19_3 , 
        \modulator_0/counter23_1 , \modulator_0/un6lto4 , 
        \modulator_0/clock_counter[2]_net_1 , 
        \modulator_0/clock_counter[3]_net_1 , 
        \modulator_0/output_signal_1_sqmuxa_0_0 , 
        \modulator_0/un6lt15 , \modulator_0/N_89 , 
        \modulator_0/clock_counter_c13 , \modulator_0/counter19 , 
        \modulator_0/clock_counter_n14 , 
        \modulator_0/clock_counter_n13 , 
        \modulator_0/clock_counter_c12 , 
        \modulator_0/clock_counter_n10 , 
        \modulator_0/clock_counter_c9 , \modulator_0/clock_counter_n9 , 
        \modulator_0/clock_counter_c8 , \modulator_0/clock_counter_n7 , 
        \modulator_0/clock_counter_c6 , 
        \modulator_0/clock_counter[7]_net_1 , 
        \modulator_0/clock_counter_n4 , \modulator_0/clock_counter_c3 , 
        \modulator_0/clock_counter_n2 , \modulator_0/clock_counter_c1 , 
        \modulator_0/clock_counter_n3 , \modulator_0/clock_counter_c2 , 
        \modulator_0/clock_counter_n5 , \modulator_0/clock_counter_c4 , 
        \modulator_0/clock_counter_n6 , \modulator_0/clock_counter_c5 , 
        \modulator_0/clock_counter_n8 , \modulator_0/clock_counter_c7 , 
        \modulator_0/clock_counter[8]_net_1 , 
        \modulator_0/clock_counter_n11 , 
        \modulator_0/clock_counter_c10 , 
        \modulator_0/clock_counter_n12 , 
        \modulator_0/clock_counter_c11 , \modulator_0/counter_n2 , 
        \modulator_0/counter_0_sqmuxa , \modulator_0/counter_n2_tz , 
        \modulator_0/counter[2]_net_1 , \modulator_0/counter_n3 , 
        \modulator_0/counter_c2 , \modulator_0/counter[3]_net_1 , 
        \modulator_0/counter_n4 , \modulator_0/counter_n4_tz , 
        \modulator_0/counter_n5 , \modulator_0/counter_45_0 , 
        \modulator_0/un6lt11 , \modulator_0/un6lt9 , 
        \modulator_0/clock_countere , \modulator_0/N_121 , 
        \modulator_0/clock_counter_n1 , 
        \modulator_0/clock_counter_n15 , \modulator_0/counter_n0 , 
        \modulator_0/counter_n1 , 
        \data_source_0/data_index_0[4]_net_1 , \data_source_0/I_12 , 
        \data_source_0/data_index_0[7]_net_1 , 
        \data_source_0/data_index_3[7] , \data_source_0/N_29 , 
        \data_source_0/counter_RNIK0AI3[1]_net_1 , 
        \data_source_0/data_index[1]_net_1 , 
        \data_source_0/data_index[0]_net_1 , 
        \data_source_0/data_index[3]_net_1 , 
        \data_source_0/DWACT_FINC_E[0] , 
        \data_source_0/data_index[8]_net_1 , 
        \data_source_0/DWACT_FINC_E[4] , 
        \data_source_0/tag_control_sig_2_0_4[15]_net_1 , 
        \data_source_0/N_1042 , 
        \data_source_0/tag_control_sig_2_0_7[11]_net_1 , 
        \data_source_0/N_994 , 
        \data_source_0/tag_control_sig_2_0_4[11]_net_1 , 
        \data_source_0/N_1001 , \data_source_0/N_1181 , 
        \data_source_0/N_1200 , \data_source_0/N_1160 , 
        \data_source_0/N_1191 , \data_source_0/N_1159 , 
        \data_source_0/N_1196 , \data_source_0/N_1162 , 
        \data_source_0/N_1187 , \data_source_0/N_1211 , 
        \data_source_0/N_1175 , \data_source_0/N_1206 , 
        \data_source_0/counter_n9_i_0 , 
        \data_source_0/counter[9]_net_1 , \data_source_0/N_38 , 
        \data_source_0/N_68 , \data_source_0/counter_n8_i_0 , 
        \data_source_0/N_34 , \data_source_0/counter_n8_i_a3_0_0 , 
        \data_source_0/N_69 , \data_source_0/N_87 , 
        \data_source_0/tag_control_sig_1_649_6 , 
        \data_source_0/tag_control_sig_1_649_1 , 
        \data_source_0/tag_control_sig_1_649_0 , 
        \data_source_0/tag_control_sig_1_649_5 , 
        \data_source_0/tag_control_sig_1_649_3 , 
        \data_source_0/data_index[6]_net_1 , 
        \data_source_0/data_index[7]_net_1 , 
        \data_source_0/data_index[2]_net_1 , 
        \data_source_0/data_index[9]_net_1 , 
        \data_source_0/output_data_1_sqmuxa_i_a3_4 , 
        \data_source_0/output_data_1_sqmuxa_i_a3_1 , 
        \data_source_0/N_90 , 
        \data_source_0/output_data_1_sqmuxa_i_a3_2 , 
        \data_source_0/counter_i_0[3] , \data_source_0/counter_i_0[2] , 
        \data_source_0/counter_i_0[4] , 
        \data_source_0/counter[8]_net_1 , 
        \data_source_0/counter_n9_i_a2_6 , 
        \data_source_0/counter_n9_i_a2_4 , 
        \data_source_0/counter[14]_net_1 , 
        \data_source_0/counter[13]_net_1 , 
        \data_source_0/counter_n9_i_a2_5 , 
        \data_source_0/counter_i_0[7] , \data_source_0/counter_i_0[6] , 
        \data_source_0/counter_n9_i_a2_2 , 
        \data_source_0/counter[5]_net_1 , 
        \data_source_0/counter[15]_net_1 , 
        \data_source_0/counter[12]_net_1 , 
        \data_source_0/counter[11]_net_1 , 
        \data_source_0/counter[10]_net_1 , 
        \data_source_0/tag_control_sig_2_0_46_tz_0 , 
        \data_source_0/N_1183 , 
        \data_source_0/tag_control_sig_2_0_a20_2_0[9] , 
        \data_source_0/N_1234 , \data_source_0/N_1144 , 
        \data_source_0/N_1148 , 
        \data_source_0/tag_control_sig_2_0_a20_0_0[17] , 
        \data_source_0/N_1145 , \data_source_0/N_1192 , 
        \data_source_0/tag_control_sig_2_0_a20_4_0[16] , 
        \data_source_0/N_1152 , 
        \data_source_0/tag_control_sig_2_0_a20_8_0[15] , 
        \data_source_0/tag_control_sig_2_0_a20_9_0[3] , 
        \data_source_0/N_1205 , \data_source_0/N_1142 , 
        \data_source_0/tag_control_sig_2_0_a20_12_0[19] , 
        \data_source_0/tag_control_sig_2_0_a20_3_0[18] , 
        \data_source_0/N_701_i , \data_source_0/N_1180 , 
        \data_source_0/tag_control_sig_2_0_a20_1_0[18] , 
        \data_source_0/N_1227 , \data_source_0/N_1232 , 
        \data_source_0/N_1186 , 
        \data_source_0/tag_control_sig_2_0_a20_3_0[6] , 
        \data_source_0/N_1140 , \data_source_0/N_1176 , 
        \data_source_0/tag_control_sig_2_0_a20_1_0[6] , 
        \data_source_0/N_1155 , \data_source_0/N_1171 , 
        \data_source_0/tag_control_sig_2_0_a20_10_0[5] , 
        \data_source_0/N_1138 , \data_source_0/N_1177 , 
        \data_source_0/tag_control_sig_2_0_a20_6_0[1] , 
        \data_source_0/N_1133 , 
        \data_source_0/tag_control_sig_2_0_a20_7_0[4] , 
        \data_source_0/tag_control_sig_2_0_a20_8_0[4] , 
        \data_source_0/N_1136 , \data_source_0/N_1134 , 
        \data_source_0/N_1139 , \data_source_0/N_1132 , 
        \data_source_0/tag_control_sig_2_0_a20_6_0[7] , 
        \data_source_0/tag_control_sig_2_0_a20_2_1[12] , 
        \data_source_0/tag_control_sig_2_0_a20_2_0[12] , 
        \data_source_0/N_1193 , 
        \data_source_0/tag_control_sig_2_0_a20_4_1[18] , 
        \data_source_0/data_index[4]_net_1 , 
        \data_source_0/tag_control_sig_2_0_a20_4_0[18] , 
        \data_source_0/tag_control_sig_2_0_a20_1_0[19] , 
        \data_source_0/N_1182 , 
        \data_source_0/tag_control_sig_2_0_12[19] , 
        \data_source_0/tag_control_sig_2_0_3[19] , 
        \data_source_0/tag_control_sig_2_0_2[19] , 
        \data_source_0/tag_control_sig_2_0_8[19] , 
        \data_source_0/tag_control_sig_2_0_11[19] , 
        \data_source_0/tag_control_sig_RNO_3[19]_net_1 , 
        \data_source_0/N_1010 , 
        \data_source_0/tag_control_sig_2_0_7[19] , 
        \data_source_0/tag_control_sig_2_0_10[19] , 
        \data_source_0/N_1056 , \data_source_0/N_883 , 
        \data_source_0/tag_control_sig_2_0_4[19] , 
        \data_source_0/N_1125 , \data_source_0/N_1117 , 
        \data_source_0/tag_control_sig_2_0_1[19] , 
        \data_source_0/N_860 , \data_source_0/N_868_1 , 
        \data_source_0/N_1120 , \data_source_0/N_1207 , 
        \data_source_0/tag_control_sig_RNO_12[19]_net_1 , 
        \data_source_0/tag_control_sig_2_0_a20_0_0[19] , 
        \data_source_0/N_1074_2 , \data_source_0/N_1129 , 
        \data_source_0/N_1237 , \data_source_0/N_1122 , 
        \data_source_0/tag_control_sig_2_0_14[18] , 
        \data_source_0/tag_control_sig_2_0_8[18] , 
        \data_source_0/tag_control_sig_2_0_7[18] , 
        \data_source_0/tag_control_sig_2_0_11[18] , 
        \data_source_0/N_1109 , \data_source_0/N_1113 , 
        \data_source_0/tag_control_sig_2_0_6[18] , 
        \data_source_0/tag_control_sig_2_0_10[18] , 
        \data_source_0/N_1111 , \data_source_0/N_1105 , 
        \data_source_0/tag_control_sig_2_0_3[18] , 
        \data_source_0/tag_control_sig_2_0_9[18] , 
        \data_source_0/N_1110 , \data_source_0/N_886 , 
        \data_source_0/tag_control_sig_2_0_2[18] , 
        \data_source_0/N_1243 , 
        \data_source_0/tag_control_sig_2_0_0[18] , 
        \data_source_0/N_1174 , \data_source_0/N_1102 , 
        \data_source_0/N_1189 , \data_source_0/N_1103 , 
        \data_source_0/N_1230 , \data_source_0/N_1114 , 
        \data_source_0/N_1188 , \data_source_0/N_1115 , 
        \data_source_0/N_1027 , 
        \data_source_0/tag_control_sig_2_0_13[16] , 
        \data_source_0/tag_control_sig_2_0_5[16] , 
        \data_source_0/tag_control_sig_2_0_4[16] , 
        \data_source_0/tag_control_sig_2_0_11[16] , 
        \data_source_0/tag_control_sig_RNO_17[16]_net_1 , 
        \data_source_0/N_1073 , 
        \data_source_0/tag_control_sig_2_0_7[16] , 
        \data_source_0/tag_control_sig_2_0_9[16] , 
        \data_source_0/N_1080 , \data_source_0/N_1083 , 
        \data_source_0/tag_control_sig_2_0_2[16] , 
        \data_source_0/tag_control_sig_2_0_8[16] , 
        \data_source_0/N_1075 , \data_source_0/N_1076 , 
        \data_source_0/tag_control_sig_2_0_1[16] , 
        \data_source_0/N_759 , \data_source_0/N_1082 , 
        \data_source_0/N_1202 , \data_source_0/N_1078 , 
        \data_source_0/N_921 , \data_source_0/N_1218 , 
        \data_source_0/N_1081 , \data_source_0/N_822 , 
        \data_source_0/N_1072 , 
        \data_source_0/tag_control_sig_2_0_a20_1_0[16] , 
        \data_source_0/N_1028 , 
        \data_source_0/tag_control_sig_2_0_15[15] , 
        \data_source_0/tag_control_sig_2_0_3[15] , 
        \data_source_0/tag_control_sig_2_0_12[15] , 
        \data_source_0/tag_control_sig_2_0_14[15] , 
        \data_source_0/tag_control_sig_2_0_0[15] , 
        \data_source_0/N_1062 , 
        \data_source_0/tag_control_sig_2_0_10[15] , 
        \data_source_0/tag_control_sig_2_0_13[15] , 
        \data_source_0/N_1064 , \data_source_0/N_1071 , 
        \data_source_0/tag_control_sig_2_0_8[15] , 
        \data_source_0/N_1061 , 
        \data_source_0/tag_control_sig_2_0_6[15] , 
        \data_source_0/N_1068 , \data_source_0/N_1057 , 
        \data_source_0/tag_control_sig_2_0_2[15] , 
        \data_source_0/N_1225 , \data_source_0/N_1063 , 
        \data_source_0/N_1059 , \data_source_0/N_1201 , 
        \data_source_0/N_1055 , \data_source_0/N_1209 , 
        \data_source_0/N_1066 , \data_source_0/N_778 , 
        \data_source_0/N_1173 , \data_source_0/N_1058 , 
        \data_source_0/tag_control_sig_2_0_12[12] , 
        \data_source_0/tag_control_sig_2_0_1[12] , 
        \data_source_0/tag_control_sig_2_0_0[12] , 
        \data_source_0/tag_control_sig_2_0_9[12] , 
        \data_source_0/tag_control_sig_2_0_11[12] , 
        \data_source_0/N_1015 , 
        \data_source_0/tag_control_sig_RNO_4[12]_net_1 , 
        \data_source_0/tag_control_sig_2_0_7[12] , 
        \data_source_0/tag_control_sig_2_0_10[12] , 
        \data_source_0/N_1018 , \data_source_0/N_1019 , 
        \data_source_0/tag_control_sig_2_0_4[12] , 
        \data_source_0/N_1006 , \data_source_0/N_1013 , 
        \data_source_0/tag_control_sig_2_0_2[12] , 
        \data_source_0/N_1014 , \data_source_0/N_873 , 
        \data_source_0/N_1213 , \data_source_0/N_1007 , 
        \data_source_0/tag_control_sig_2_0_a20_1_1[12] , 
        \data_source_0/tag_control_sig_2_0_a20_1_0[12] , 
        \data_source_0/N_835 , 
        \data_source_0/tag_control_sig_2_0_12[10] , 
        \data_source_0/tag_control_sig_2_0_6[10] , 
        \data_source_0/tag_control_sig_2_0_5[10] , 
        \data_source_0/tag_control_sig_2_0_9[10] , 
        \data_source_0/N_978 , \data_source_0/N_979 , 
        \data_source_0/tag_control_sig_2_0_4[10] , 
        \data_source_0/tag_control_sig_2_0_8[10] , 
        \data_source_0/N_980 , \data_source_0/N_976 , 
        \data_source_0/tag_control_sig_2_0_2[10] , 
        \data_source_0/tag_control_sig_2_0_7[10] , 
        \data_source_0/N_779 , \data_source_0/N_1204 , 
        \data_source_0/tag_control_sig_2_0_0[10] , 
        \data_source_0/N_726 , \data_source_0/N_982 , 
        \data_source_0/N_1195 , \data_source_0/N_1163 , 
        \data_source_0/N_975 , \data_source_0/N_1220 , 
        \data_source_0/N_1219 , \data_source_0/N_985 , 
        \data_source_0/N_984 , 
        \data_source_0/tag_control_sig_2_0_a20_3_1[10] , 
        \data_source_0/tag_control_sig_2_0_a20_3_0[10] , 
        \data_source_0/N_981 , 
        \data_source_0/tag_control_sig_2_0_13[8] , 
        \data_source_0/tag_control_sig_2_0_5[8] , 
        \data_source_0/tag_control_sig_2_0_4[8] , 
        \data_source_0/tag_control_sig_2_0_11[8] , 
        \data_source_0/N_950 , \data_source_0/N_951 , 
        \data_source_0/tag_control_sig_2_0_7[8] , 
        \data_source_0/tag_control_sig_2_0_9[8] , 
        \data_source_0/N_945 , \data_source_0/N_879 , 
        \data_source_0/tag_control_sig_2_0_3[8] , 
        \data_source_0/tag_control_sig_2_0_8[8] , 
        \data_source_0/N_955 , \data_source_0/N_953 , 
        \data_source_0/tag_control_sig_2_0_1[8] , 
        \data_source_0/N_943 , \data_source_0/N_729 , 
        \data_source_0/N_949 , \data_source_0/N_947 , 
        \data_source_0/N_800 , \data_source_0/N_954 , 
        \data_source_0/N_785 , \data_source_0/N_1199 , 
        \data_source_0/N_952 , 
        \data_source_0/tag_control_sig_2_0_12[7] , 
        \data_source_0/tag_control_sig_2_0_6[7] , 
        \data_source_0/tag_control_sig_2_0_5[7] , 
        \data_source_0/tag_control_sig_2_0_9[7] , 
        \data_source_0/tag_control_sig_2_0_11[7] , 
        \data_source_0/tag_control_sig_2_0_0[7] , 
        \data_source_0/N_936 , 
        \data_source_0/tag_control_sig_2_0_8[7] , 
        \data_source_0/N_939 , \data_source_0/N_927 , 
        \data_source_0/tag_control_sig_2_0_4[7] , 
        \data_source_0/N_930 , \data_source_0/N_929 , 
        \data_source_0/tag_control_sig_2_0_1[7] , 
        \data_source_0/N_935 , \data_source_0/N_766 , 
        \data_source_0/N_931 , 
        \data_source_0/tag_control_sig_2_0_a20_4_1[7] , 
        \data_source_0/tag_control_sig_2_0_a20_4_0[7] , 
        \data_source_0/N_938 , \data_source_0/N_1179 , 
        \data_source_0/N_819 , \data_source_0/N_1161 , 
        \data_source_0/tag_control_sig_2_0_2_tz[7] , 
        \data_source_0/N_941 , 
        \data_source_0/tag_control_sig_2_0_15[6] , 
        \data_source_0/tag_control_sig_2_0_9[6] , 
        \data_source_0/tag_control_sig_2_0_8[6] , 
        \data_source_0/tag_control_sig_2_0_12[6] , 
        \data_source_0/N_833 , 
        \data_source_0/tag_control_sig_2_0_6[6] , 
        \data_source_0/tag_control_sig_2_0_11[6] , 
        \data_source_0/N_856 , \data_source_0/N_920 , 
        \data_source_0/tag_control_sig_2_0_5[6] , 
        \data_source_0/tag_control_sig_2_0_10[6] , 
        \data_source_0/N_915 , \data_source_0/N_914 , 
        \data_source_0/tag_control_sig_2_0_3[6] , 
        \data_source_0/N_817 , \data_source_0/N_903 , 
        \data_source_0/tag_control_sig_2_0_0[6] , 
        \data_source_0/N_1197 , \data_source_0/N_923 , 
        \data_source_0/N_1242 , \data_source_0/N_925 , 
        \data_source_0/N_1233 , \data_source_0/N_919 , 
        \data_source_0/N_917 , \data_source_0/N_924 , 
        \data_source_0/tag_control_sig_2_0_13[5] , 
        \data_source_0/tag_control_sig_2_0_4[5] , 
        \data_source_0/tag_control_sig_2_0_3[5] , 
        \data_source_0/tag_control_sig_2_0_9[5] , 
        \data_source_0/tag_control_sig_2_0_12[5] , 
        \data_source_0/tag_control_sig_2_0_0[5] , 
        \data_source_0/N_910 , 
        \data_source_0/tag_control_sig_2_0_7[5] , 
        \data_source_0/tag_control_sig_2_0_11[5] , 
        \data_source_0/N_907 , \data_source_0/N_909 , 
        \data_source_0/tag_control_sig_2_0_6[5] , 
        \data_source_0/N_897 , \data_source_0/N_908 , 
        \data_source_0/tag_control_sig_2_0_1[5] , 
        \data_source_0/tag_control_sig_2_0_a20_3_0[5] , 
        \data_source_0/N_901_1 , \data_source_0/N_911 , 
        \data_source_0/N_904 , \data_source_0/N_804 , 
        \data_source_0/N_902 , 
        \data_source_0/tag_control_sig_2_0_a20_1_1[5] , 
        \data_source_0/tag_control_sig_2_0_a20_1_0[5] , 
        \data_source_0/N_900 , 
        \data_source_0/tag_control_sig_2_0_13[4] , 
        \data_source_0/tag_control_sig_2_0_5[4] , 
        \data_source_0/tag_control_sig_2_0_4[4] , 
        \data_source_0/tag_control_sig_2_0_11[4] , 
        \data_source_0/N_889 , \data_source_0/N_895 , 
        \data_source_0/tag_control_sig_2_0_7[4] , 
        \data_source_0/tag_control_sig_2_0_9[4] , 
        \data_source_0/N_887 , 
        \data_source_0/tag_control_sig_2_0_3[4] , 
        \data_source_0/tag_control_sig_2_0_8[4] , 
        \data_source_0/N_881 , \data_source_0/N_764 , 
        \data_source_0/tag_control_sig_2_0_0[4] , 
        \data_source_0/N_894 , \data_source_0/N_888 , 
        \data_source_0/tag_control_sig_RNO_11[4]_net_1 , 
        \data_source_0/N_783 , \data_source_0/N_996_1 , 
        \data_source_0/tag_control_sig_2_0_13[2] , 
        \data_source_0/tag_control_sig_2_0_2[2] , 
        \data_source_0/tag_control_sig_2_0_1[2] , 
        \data_source_0/tag_control_sig_2_0_10[2] , 
        \data_source_0/tag_control_sig_2_0_12[2] , 
        \data_source_0/tag_control_sig_2_0_0[2] , 
        \data_source_0/N_859 , 
        \data_source_0/tag_control_sig_2_0_7[2] , 
        \data_source_0/tag_control_sig_2_0_11[2] , 
        \data_source_0/N_863 , \data_source_0/N_862 , 
        \data_source_0/tag_control_sig_2_0_6[2] , 
        \data_source_0/tag_control_sig_RNO_13[2]_net_1 , 
        \data_source_0/N_851 , 
        \data_source_0/tag_control_sig_2_0_3[2] , 
        \data_source_0/N_1190 , \data_source_0/N_832 , 
        \data_source_0/tag_control_sig_2_0_a20_3_0[2] , 
        \data_source_0/N_853_2 , \data_source_0/N_854 , 
        \data_source_0/N_849 , 
        \data_source_0/tag_control_sig_2_0_16[1] , 
        \data_source_0/tag_control_sig_2_0_10[1] , 
        \data_source_0/tag_control_sig_2_0_9[1] , 
        \data_source_0/tag_control_sig_2_0_13[1] , 
        \data_source_0/N_848 , \data_source_0/N_847 , 
        \data_source_0/tag_control_sig_2_0_7[1] , 
        \data_source_0/tag_control_sig_2_0_12[1] , 
        \data_source_0/N_844 , \data_source_0/N_843 , 
        \data_source_0/tag_control_sig_2_0_5[1] , 
        \data_source_0/tag_control_sig_2_0_11[1] , 
        \data_source_0/tag_control_sig_2_0_3[1] , 
        \data_source_0/N_831 , 
        \data_source_0/tag_control_sig_2_0_4[1] , 
        \data_source_0/N_834 , 
        \data_source_0/tag_control_sig_2_0_2[1] , 
        \data_source_0/N_830 , \data_source_0/N_829 , 
        \data_source_0/N_1184 , \data_source_0/N_846 , 
        \data_source_0/N_1198 , \data_source_0/N_841 , 
        \data_source_0/N_837 , 
        \data_source_0/tag_control_sig_2_0_a20_2_0[19] , 
        \data_source_0/N_1135 , 
        \data_source_0/tag_control_sig_2_0_a20_2_1[18] , 
        \data_source_0/N_704_i , 
        \data_source_0/tag_control_sig_2_0_a20_2_0[18] , 
        \data_source_0/tag_control_sig_2_0_a20_2[16] , 
        \data_source_0/N_1157 , \data_source_0/data_index[5]_net_1 , 
        \data_source_0/tag_control_sig_2_0_a20_3_0[9] , 
        \data_source_0/N_1143 , 
        \data_source_0/tag_control_sig_2_0_a20_0_1[15] , 
        \data_source_0/N_707_i , 
        \data_source_0/tag_control_sig_2_0_a20_5_0[10] , 
        \data_source_0/N_1231 , 
        \data_source_0/tag_control_sig_2_0_a20_4_0[10] , 
        \data_source_0/N_1239 , \data_source_0/N_703_i , 
        \data_source_0/tag_control_sig_2_0_a20_10_0[8] , 
        \data_source_0/N_1156 , \data_source_0/N_1141 , 
        \data_source_0/tag_control_sig_2_0_a20_6_0[8] , 
        \data_source_0/tag_control_sig_2_0_a20_4_0[8] , 
        \data_source_0/N_1208 , \data_source_0/N_1238 , 
        \data_source_0/tag_control_sig_2_0_a20_3_0[7] , 
        \data_source_0/tag_control_sig_2_0_a20_2_0[7] , 
        \data_source_0/tag_control_sig_2_0_a20_0[7] , 
        \data_source_0/tag_control_sig_2_0_a20_2_0[6] , 
        \data_source_0/N_1137 , 
        \data_source_0/tag_control_sig_2_0_14[17] , 
        \data_source_0/tag_control_sig_2_0_8[17] , 
        \data_source_0/tag_control_sig_2_0_7[17] , 
        \data_source_0/tag_control_sig_2_0_11[17] , 
        \data_source_0/N_1096 , \data_source_0/N_1094 , 
        \data_source_0/tag_control_sig_2_0_5[17] , 
        \data_source_0/tag_control_sig_2_0_10[17] , 
        \data_source_0/N_1088 , \data_source_0/N_1089 , 
        \data_source_0/tag_control_sig_2_0_3[17] , 
        \data_source_0/tag_control_sig_2_0_9[17] , 
        \data_source_0/N_1091 , \data_source_0/N_1090 , 
        \data_source_0/tag_control_sig_2_0_2[17] , 
        \data_source_0/N_1100 , \data_source_0/N_1099 , 
        \data_source_0/N_1098 , \data_source_0/N_1097 , 
        \data_source_0/N_1101 , \data_source_0/N_748 , 
        \data_source_0/N_1086 , \data_source_0/N_1092 , 
        \data_source_0/tag_control_sig_2_0_14[14] , 
        \data_source_0/tag_control_sig_2_0_5[14] , 
        \data_source_0/tag_control_sig_2_0_4[14] , 
        \data_source_0/tag_control_sig_2_0_10[14] , 
        \data_source_0/tag_control_sig_2_0_13[14] , 
        \data_source_0/tag_control_sig_2_0_1[14] , 
        \data_source_0/tag_control_sig_2_0_0[14] , 
        \data_source_0/tag_control_sig_2_0_8[14] , 
        \data_source_0/tag_control_sig_2_0_12[14] , 
        \data_source_0/N_1044 , \data_source_0/N_1041 , 
        \data_source_0/tag_control_sig_2_0_6[14] , 
        \data_source_0/N_1040 , \data_source_0/N_1049 , 
        \data_source_0/tag_control_sig_2_0_3[14] , 
        \data_source_0/N_1046 , \data_source_0/N_802 , 
        \data_source_0/N_1052 , \data_source_0/N_1050 , 
        \data_source_0/N_1045 , \data_source_0/N_1215 , 
        \data_source_0/N_1038 , 
        \data_source_0/tag_control_sig_2_0_16[13] , 
        \data_source_0/tag_control_sig_2_0_7[13] , 
        \data_source_0/tag_control_sig_2_0_6[13] , 
        \data_source_0/tag_control_sig_2_0_12[13] , 
        \data_source_0/tag_control_sig_2_0_15[13] , 
        \data_source_0/tag_control_sig_2_0_3[13] , 
        \data_source_0/tag_control_sig_2_0_2[13] , 
        \data_source_0/tag_control_sig_2_0_10[13] , 
        \data_source_0/tag_control_sig_2_0_14[13] , 
        \data_source_0/N_1030 , \data_source_0/N_1033 , 
        \data_source_0/tag_control_sig_2_0_9[13] , 
        \data_source_0/N_1026 , 
        \data_source_0/tag_control_sig_2_0_5[13] , 
        \data_source_0/N_1035 , \data_source_0/N_1025 , 
        \data_source_0/tag_control_sig_2_0_1[13] , 
        \data_source_0/N_1024 , \data_source_0/N_1031 , 
        \data_source_0/N_1235 , \data_source_0/N_1023 , 
        \data_source_0/N_1034 , \data_source_0/N_1223 , 
        \data_source_0/N_1224 , \data_source_0/N_1020 , 
        \data_source_0/N_1021 , 
        \data_source_0/tag_control_sig_2_0_17[11] , 
        \data_source_0/tag_control_sig_2_0_6[11] , 
        \data_source_0/tag_control_sig_2_0_5[11] , 
        \data_source_0/tag_control_sig_2_0_14[11] , 
        \data_source_0/tag_control_sig_2_0_16[11] , 
        \data_source_0/tag_control_sig_2_0_2[11] , 
        \data_source_0/tag_control_sig_2_0_1[11] , 
        \data_source_0/tag_control_sig_2_0_12[11] , 
        \data_source_0/tag_control_sig_2_0_15[11] , 
        \data_source_0/tag_control_sig_2_0_0[11] , 
        \data_source_0/N_991 , 
        \data_source_0/tag_control_sig_2_0_9[11] , 
        \data_source_0/N_990 , \data_source_0/N_997 , 
        \data_source_0/N_988 , \data_source_0/N_987 , 
        \data_source_0/N_993 , \data_source_0/N_1000 , 
        \data_source_0/N_872 , \data_source_0/N_1185 , 
        \data_source_0/N_995 , \data_source_0/N_1005 , 
        \data_source_0/tag_control_sig_2_0_14[9] , 
        \data_source_0/tag_control_sig_2_0_3[9] , 
        \data_source_0/tag_control_sig_2_0_2[9] , 
        \data_source_0/tag_control_sig_2_0_11[9] , 
        \data_source_0/tag_control_sig_2_0_13[9] , 
        \data_source_0/tag_control_sig_2_0_1[9] , 
        \data_source_0/tag_control_sig_2_0_0[9] , 
        \data_source_0/tag_control_sig_2_0_8[9] , 
        \data_source_0/tag_control_sig_2_0_12[9] , 
        \data_source_0/N_962 , \data_source_0/N_969 , 
        \data_source_0/tag_control_sig_2_0_7[9] , 
        \data_source_0/N_968 , \data_source_0/N_967 , 
        \data_source_0/tag_control_sig_2_0_5[9] , 
        \data_source_0/N_1229 , \data_source_0/N_1178 , 
        \data_source_0/N_960 , \data_source_0/N_961 , 
        \data_source_0/N_970 , \data_source_0/N_965 , 
        \data_source_0/N_777 , \data_source_0/N_957 , 
        \data_source_0/N_1245 , \data_source_0/N_816 , 
        \data_source_0/N_964 , 
        \data_source_0/tag_control_sig_2_0_14[3] , 
        \data_source_0/tag_control_sig_2_0_8[3] , 
        \data_source_0/tag_control_sig_2_0_7[3] , 
        \data_source_0/tag_control_sig_2_0_11[3] , 
        \data_source_0/N_875 , 
        \data_source_0/tag_control_sig_2_0_5[3] , 
        \data_source_0/tag_control_sig_2_0_10[3] , 
        \data_source_0/N_867 , \data_source_0/N_876 , 
        \data_source_0/tag_control_sig_2_0_3[3] , 
        \data_source_0/tag_control_sig_2_0_9[3] , 
        \data_source_0/tag_control_sig_2_0_1[3] , 
        \data_source_0/N_757 , 
        \data_source_0/tag_control_sig_2_0_0[3] , 
        \data_source_0/N_869 , \data_source_0/N_868 , 
        \data_source_0/N_877 , \data_source_0/N_808 , 
        \data_source_0/N_865 , \data_source_0/N_1240 , 
        \data_source_0/N_870 , 
        \data_source_0/tag_control_sig_2_0_14[0] , 
        \data_source_0/tag_control_sig_2_0_10[0] , 
        \data_source_0/tag_control_sig_2_0_11[0] , 
        \data_source_0/tag_control_sig_2_0_13[0] , 
        \data_source_0/tag_control_sig_2_0_1[0] , 
        \data_source_0/tag_control_sig_2_0_0[0] , 
        \data_source_0/tag_control_sig_2_0_8[0] , 
        \data_source_0/tag_control_sig_2_0_12[0] , 
        \data_source_0/N_811 , \data_source_0/N_825 , 
        \data_source_0/tag_control_sig_2_0_7[0] , 
        \data_source_0/N_827 , 
        \data_source_0/tag_control_sig_2_0_6[0] , 
        \data_source_0/tag_control_sig_2_0_5[0] , 
        \data_source_0/N_815 , \data_source_0/N_823 , 
        \data_source_0/tag_control_sig_2_0_3[0] , 
        \data_source_0/N_813 , \data_source_0/N_818 , 
        \data_source_0/N_1244 , \data_source_0/N_820 , 
        \data_source_0/tag_control_sig_2_0_a20_3_2[9] , 
        \data_source_0/tag_control_sig_2_0_a20_3_0[3] , 
        \data_source_0/tag_control_sig_2_0_a20_2_0[3] , 
        \data_source_0/tag_control_sig_2_0_a20_0[0] , 
        \data_source_0/tag_control_sig_2_0_a20_4_1[17] , 
        \data_source_0/tag_control_sig_2_0_a20_2_1[17] , 
        \data_source_0/tag_control_sig_2_0_a20_9_2[16] , 
        \data_source_0/N_1149 , \data_source_0/N_18 , 
        \data_source_0/N_53_i , \data_source_0/N_73 , 
        \data_source_0/N_12 , \data_source_0/N_10 , 
        \data_source_0/N_39 , \data_source_0/N_813_1 , 
        \data_source_0/N_919_1 , \data_source_0/N_1040_1 , 
        \data_source_0/tag_control_sig_2[0] , 
        \data_source_0/tag_control_sig_2[3] , 
        \data_source_0/tag_control_sig_2[9] , 
        \data_source_0/tag_control_sig_2[11] , 
        \data_source_0/tag_control_sig_2[13] , 
        \data_source_0/tag_control_sig_2[14] , \data_source_0/N_668 , 
        \data_source_0/tag_control_sig_2[1] , 
        \data_source_0/tag_control_sig_2[2] , 
        \data_source_0/tag_control_sig_2[4] , 
        \data_source_0/tag_control_sig_2[5] , 
        \data_source_0/tag_control_sig_2[6] , 
        \data_source_0/tag_control_sig_2[7] , 
        \data_source_0/tag_control_sig_2[8] , 
        \data_source_0/tag_control_sig_2[10] , 
        \data_source_0/tag_control_sig_2[12] , 
        \data_source_0/tag_control_sig_2[15] , 
        \data_source_0/tag_control_sig_2[16] , 
        \data_source_0/tag_control_sig_2[17] , 
        \data_source_0/tag_control_sig_2[18] , 
        \data_source_0/tag_control_sig_2[19] , \data_source_0/N_807 , 
        \data_source_0/N_1151 , \data_source_0/N_1154 , 
        \data_source_0/N_1217 , \data_source_0/N_771 , 
        \data_source_0/tag_control_sig_1_3[649] , \data_source_0/N_26 , 
        \data_source_0/counter_i_0[0] , \data_source_0/counter_i_0[1] , 
        \data_source_0/N_24 , \data_source_0/N_31 , 
        \data_source_0/N_22 , \data_source_0/N_32 , 
        \data_source_0/N_20 , \data_source_0/N_33 , 
        \data_source_0/N_16 , \data_source_0/N_35 , 
        \data_source_0/N_14 , \data_source_0/N_36 , 
        \data_source_0/N_1210 , 
        \data_source_0/tag_control_sig_2_0_a20_9_0[1] , 
        \data_source_0/tag_control_sig_2_0_a20_10_0[1] , 
        \data_source_0/N_534_tz , \data_source_0/N_1226 , 
        \data_source_0/N_1123_1 , \data_source_0/counter_n15 , 
        \data_source_0/N_44 , \data_source_0/counter_n14 , 
        \data_source_0/N_43 , \data_source_0/counter_n13 , 
        \data_source_0/N_42 , \data_source_0/counter_n12 , 
        \data_source_0/N_41 , \data_source_0/counter_n11 , 
        \data_source_0/N_40 , \data_source_0/counter_n10 , 
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 , 
        \data_source_0/data_index_3[1] , \data_source_0/I_5 , 
        \data_source_0/data_index_3[3] , \data_source_0/I_9 , 
        \data_source_0/I_20 , \data_source_0/data_index_3[9] , 
        \data_source_0/I_26 , \data_source_0/tag_data_buf_1_4[1] , 
        \data_source_0/tag_data_buf_1[0]_net_1 , 
        \data_source_0/tag_data_buf_1_4[2] , 
        \data_source_0/tag_data_buf_1[1]_net_1 , 
        \data_source_0/tag_data_buf_1_4[3] , 
        \data_source_0/tag_data_buf_1[2]_net_1 , 
        \data_source_0/tag_data_buf_1_4[4] , 
        \data_source_0/tag_data_buf_1[3]_net_1 , 
        \data_source_0/tag_data_buf_1_4[5] , 
        \data_source_0/tag_data_buf_1[4]_net_1 , 
        \data_source_0/tag_data_buf_1_4[6] , 
        \data_source_0/tag_data_buf_1[5]_net_1 , 
        \data_source_0/tag_data_buf_1_4[7] , 
        \data_source_0/tag_data_buf_1[6]_net_1 , 
        \data_source_0/tag_data_buf_2_4[1] , 
        \data_source_0/tag_data_buf_2[0]_net_1 , 
        \data_source_0/tag_data_buf_2_4[2] , 
        \data_source_0/tag_data_buf_2[1]_net_1 , 
        \data_source_0/tag_data_buf_2_4[3] , 
        \data_source_0/tag_data_buf_2[2]_net_1 , 
        \data_source_0/tag_data_buf_2_4[4] , 
        \data_source_0/tag_data_buf_2[3]_net_1 , 
        \data_source_0/tag_data_buf_2_4[5] , 
        \data_source_0/tag_data_buf_2[4]_net_1 , 
        \data_source_0/tag_data_buf_2_4[6] , 
        \data_source_0/tag_data_buf_2[5]_net_1 , 
        \data_source_0/tag_data_buf_2_4[7] , 
        \data_source_0/tag_data_buf_2[6]_net_1 , 
        \data_source_0/tag_data_buf_3_4[1] , 
        \data_source_0/tag_data_buf_3[0]_net_1 , 
        \data_source_0/tag_data_buf_3_4[2] , 
        \data_source_0/tag_data_buf_3[1]_net_1 , 
        \data_source_0/tag_data_buf_3_4[3] , 
        \data_source_0/tag_data_buf_3[2]_net_1 , 
        \data_source_0/tag_data_buf_3_4[4] , 
        \data_source_0/tag_data_buf_3[3]_net_1 , 
        \data_source_0/tag_data_buf_3_4[5] , 
        \data_source_0/tag_data_buf_3[4]_net_1 , 
        \data_source_0/tag_data_buf_3_4[6] , 
        \data_source_0/tag_data_buf_3[5]_net_1 , 
        \data_source_0/tag_data_buf_3_4[7] , 
        \data_source_0/tag_data_buf_3[6]_net_1 , 
        \data_source_0/tag_data_buf_4_4[1] , 
        \data_source_0/tag_data_buf_4[0]_net_1 , 
        \data_source_0/tag_data_buf_4_4[2] , 
        \data_source_0/tag_data_buf_4[1]_net_1 , 
        \data_source_0/tag_data_buf_4_4[3] , 
        \data_source_0/tag_data_buf_4[2]_net_1 , 
        \data_source_0/tag_data_buf_4_4[4] , 
        \data_source_0/tag_data_buf_4[3]_net_1 , 
        \data_source_0/tag_data_buf_4_4[5] , 
        \data_source_0/tag_data_buf_4[4]_net_1 , 
        \data_source_0/tag_data_buf_4_4[6] , 
        \data_source_0/tag_data_buf_4[5]_net_1 , 
        \data_source_0/tag_data_buf_4_4[7] , 
        \data_source_0/tag_data_buf_4[6]_net_1 , 
        \data_source_0/tag_data_buf_5_4[1] , 
        \data_source_0/tag_data_buf_5[0]_net_1 , 
        \data_source_0/tag_data_buf_5_4[2] , 
        \data_source_0/tag_data_buf_5[1]_net_1 , 
        \data_source_0/tag_data_buf_5_4[3] , 
        \data_source_0/tag_data_buf_5[2]_net_1 , 
        \data_source_0/tag_data_buf_5_4[4] , 
        \data_source_0/tag_data_buf_5[3]_net_1 , 
        \data_source_0/tag_data_buf_5_4[5] , 
        \data_source_0/tag_data_buf_5[4]_net_1 , 
        \data_source_0/tag_data_buf_5_4[6] , 
        \data_source_0/tag_data_buf_5[5]_net_1 , 
        \data_source_0/tag_data_buf_5_4[7] , 
        \data_source_0/tag_data_buf_5[6]_net_1 , 
        \data_source_0/tag_data_buf_6_4[1] , 
        \data_source_0/tag_data_buf_6[0]_net_1 , 
        \data_source_0/tag_data_buf_6_4[2] , 
        \data_source_0/tag_data_buf_6[1]_net_1 , 
        \data_source_0/tag_data_buf_6_4[3] , 
        \data_source_0/tag_data_buf_6[2]_net_1 , 
        \data_source_0/tag_data_buf_6_4[4] , 
        \data_source_0/tag_data_buf_6[3]_net_1 , 
        \data_source_0/tag_data_buf_6_4[5] , 
        \data_source_0/tag_data_buf_6[4]_net_1 , 
        \data_source_0/tag_data_buf_6_4[6] , 
        \data_source_0/tag_data_buf_6[5]_net_1 , 
        \data_source_0/tag_data_buf_6_4[7] , 
        \data_source_0/tag_data_buf_6[6]_net_1 , 
        \data_source_0/tag_data_buf_7_4[1] , 
        \data_source_0/tag_data_buf_7[0]_net_1 , 
        \data_source_0/tag_data_buf_7_4[2] , 
        \data_source_0/tag_data_buf_7[1]_net_1 , 
        \data_source_0/tag_data_buf_7_4[3] , 
        \data_source_0/tag_data_buf_7[2]_net_1 , 
        \data_source_0/tag_data_buf_7_4[4] , 
        \data_source_0/tag_data_buf_7[3]_net_1 , 
        \data_source_0/tag_data_buf_7_4[5] , 
        \data_source_0/tag_data_buf_7[4]_net_1 , 
        \data_source_0/tag_data_buf_7_4[6] , 
        \data_source_0/tag_data_buf_7[5]_net_1 , 
        \data_source_0/tag_data_buf_7_4[7] , 
        \data_source_0/tag_data_buf_7[6]_net_1 , 
        \data_source_0/tag_data_buf_8_4[1] , 
        \data_source_0/tag_data_buf_8[0]_net_1 , 
        \data_source_0/tag_data_buf_8_4[2] , 
        \data_source_0/tag_data_buf_8[1]_net_1 , 
        \data_source_0/tag_data_buf_8_4[3] , 
        \data_source_0/tag_data_buf_8[2]_net_1 , 
        \data_source_0/tag_data_buf_8_4[4] , 
        \data_source_0/tag_data_buf_8[3]_net_1 , 
        \data_source_0/tag_data_buf_8_4[5] , 
        \data_source_0/tag_data_buf_8[4]_net_1 , 
        \data_source_0/tag_data_buf_8_4[6] , 
        \data_source_0/tag_data_buf_8[5]_net_1 , 
        \data_source_0/tag_data_buf_8_4[7] , 
        \data_source_0/tag_data_buf_8[6]_net_1 , 
        \data_source_0/tag_data_buf_10_4[1] , 
        \data_source_0/tag_data_buf_10[0]_net_1 , 
        \data_source_0/tag_data_buf_10_4[2] , 
        \data_source_0/tag_data_buf_10[1]_net_1 , 
        \data_source_0/tag_data_buf_10_4[3] , 
        \data_source_0/tag_data_buf_10[2]_net_1 , 
        \data_source_0/tag_data_buf_10_4[4] , 
        \data_source_0/tag_data_buf_10[3]_net_1 , 
        \data_source_0/tag_data_buf_10_4[5] , 
        \data_source_0/tag_data_buf_10[4]_net_1 , 
        \data_source_0/tag_data_buf_10_4[6] , 
        \data_source_0/tag_data_buf_10[5]_net_1 , 
        \data_source_0/tag_data_buf_10_4[7] , 
        \data_source_0/tag_data_buf_10[6]_net_1 , 
        \data_source_0/tag_data_buf_11_4[1] , 
        \data_source_0/tag_data_buf_11[0]_net_1 , 
        \data_source_0/tag_data_buf_11_4[2] , 
        \data_source_0/tag_data_buf_11[1]_net_1 , 
        \data_source_0/tag_data_buf_11_4[3] , 
        \data_source_0/tag_data_buf_11[2]_net_1 , 
        \data_source_0/tag_data_buf_11_4[4] , 
        \data_source_0/tag_data_buf_11[3]_net_1 , 
        \data_source_0/tag_data_buf_11_4[5] , 
        \data_source_0/tag_data_buf_11[4]_net_1 , 
        \data_source_0/tag_data_buf_11_4[6] , 
        \data_source_0/tag_data_buf_11[5]_net_1 , 
        \data_source_0/tag_data_buf_11_4[7] , 
        \data_source_0/tag_data_buf_11[6]_net_1 , 
        \data_source_0/tag_data_buf_12_4[1] , 
        \data_source_0/tag_data_buf_12[0]_net_1 , 
        \data_source_0/tag_data_buf_12_4[2] , 
        \data_source_0/tag_data_buf_12[1]_net_1 , 
        \data_source_0/tag_data_buf_12_4[3] , 
        \data_source_0/tag_data_buf_12[2]_net_1 , 
        \data_source_0/tag_data_buf_12_4[4] , 
        \data_source_0/tag_data_buf_12[3]_net_1 , 
        \data_source_0/tag_data_buf_12_4[5] , 
        \data_source_0/tag_data_buf_12[4]_net_1 , 
        \data_source_0/tag_data_buf_12_4[6] , 
        \data_source_0/tag_data_buf_12[5]_net_1 , 
        \data_source_0/tag_data_buf_12_4[7] , 
        \data_source_0/tag_data_buf_12[6]_net_1 , 
        \data_source_0/tag_data_buf_13_4[1] , 
        \data_source_0/tag_data_buf_13[0]_net_1 , 
        \data_source_0/tag_data_buf_13_4[2] , 
        \data_source_0/tag_data_buf_13[1]_net_1 , 
        \data_source_0/tag_data_buf_13_4[3] , 
        \data_source_0/tag_data_buf_13[2]_net_1 , 
        \data_source_0/tag_data_buf_13_4[4] , 
        \data_source_0/tag_data_buf_13[3]_net_1 , 
        \data_source_0/tag_data_buf_13_4[5] , 
        \data_source_0/tag_data_buf_13[4]_net_1 , 
        \data_source_0/tag_data_buf_13_4[6] , 
        \data_source_0/tag_data_buf_13[5]_net_1 , 
        \data_source_0/tag_data_buf_13_4[7] , 
        \data_source_0/tag_data_buf_13[6]_net_1 , 
        \data_source_0/tag_data_buf_14_4[1] , 
        \data_source_0/tag_data_buf_14[0]_net_1 , 
        \data_source_0/tag_data_buf_14_4[2] , 
        \data_source_0/tag_data_buf_14[1]_net_1 , 
        \data_source_0/tag_data_buf_14_4[3] , 
        \data_source_0/tag_data_buf_14[2]_net_1 , 
        \data_source_0/tag_data_buf_14_4[4] , 
        \data_source_0/tag_data_buf_14[3]_net_1 , 
        \data_source_0/tag_data_buf_14_4[5] , 
        \data_source_0/tag_data_buf_14[4]_net_1 , 
        \data_source_0/tag_data_buf_14_4[6] , 
        \data_source_0/tag_data_buf_14[5]_net_1 , 
        \data_source_0/tag_data_buf_14_4[7] , 
        \data_source_0/tag_data_buf_14[6]_net_1 , 
        \data_source_0/tag_data_buf_15_4[1] , 
        \data_source_0/tag_data_buf_15[0]_net_1 , 
        \data_source_0/tag_data_buf_15_4[2] , 
        \data_source_0/tag_data_buf_15[1]_net_1 , 
        \data_source_0/tag_data_buf_15_4[3] , 
        \data_source_0/tag_data_buf_15[2]_net_1 , 
        \data_source_0/tag_data_buf_15_4[4] , 
        \data_source_0/tag_data_buf_15[3]_net_1 , 
        \data_source_0/tag_data_buf_15_4[5] , 
        \data_source_0/tag_data_buf_15[4]_net_1 , 
        \data_source_0/tag_data_buf_15_4[6] , 
        \data_source_0/tag_data_buf_15[5]_net_1 , 
        \data_source_0/tag_data_buf_15_4[7] , 
        \data_source_0/tag_data_buf_15[6]_net_1 , 
        \data_source_0/tag_data_buf_16_4[1] , 
        \data_source_0/tag_data_buf_16[0]_net_1 , 
        \data_source_0/tag_data_buf_16_4[2] , 
        \data_source_0/tag_data_buf_16[1]_net_1 , 
        \data_source_0/tag_data_buf_16_4[3] , 
        \data_source_0/tag_data_buf_16[2]_net_1 , 
        \data_source_0/tag_data_buf_16_4[4] , 
        \data_source_0/tag_data_buf_16[3]_net_1 , 
        \data_source_0/tag_data_buf_16_4[5] , 
        \data_source_0/tag_data_buf_16[4]_net_1 , 
        \data_source_0/tag_data_buf_16_4[6] , 
        \data_source_0/tag_data_buf_16[5]_net_1 , 
        \data_source_0/tag_data_buf_16_4[7] , 
        \data_source_0/tag_data_buf_16[6]_net_1 , 
        \data_source_0/tag_data_buf_17_4[1] , 
        \data_source_0/tag_data_buf_17[0]_net_1 , 
        \data_source_0/tag_data_buf_17_4[2] , 
        \data_source_0/tag_data_buf_17[1]_net_1 , 
        \data_source_0/tag_data_buf_17_4[3] , 
        \data_source_0/tag_data_buf_17[2]_net_1 , 
        \data_source_0/tag_data_buf_17_4[4] , 
        \data_source_0/tag_data_buf_17[3]_net_1 , 
        \data_source_0/tag_data_buf_17_4[5] , 
        \data_source_0/tag_data_buf_17[4]_net_1 , 
        \data_source_0/tag_data_buf_17_4[6] , 
        \data_source_0/tag_data_buf_17[5]_net_1 , 
        \data_source_0/tag_data_buf_17_4[7] , 
        \data_source_0/tag_data_buf_17[6]_net_1 , 
        \data_source_0/tag_data_buf_18_4[1] , 
        \data_source_0/tag_data_buf_18[0]_net_1 , 
        \data_source_0/tag_data_buf_18_4[2] , 
        \data_source_0/tag_data_buf_18[1]_net_1 , 
        \data_source_0/tag_data_buf_18_4[3] , 
        \data_source_0/tag_data_buf_18[2]_net_1 , 
        \data_source_0/tag_data_buf_18_4[4] , 
        \data_source_0/tag_data_buf_18[3]_net_1 , 
        \data_source_0/tag_data_buf_18_4[5] , 
        \data_source_0/tag_data_buf_18[4]_net_1 , 
        \data_source_0/tag_data_buf_18_4[6] , 
        \data_source_0/tag_data_buf_18[5]_net_1 , 
        \data_source_0/tag_data_buf_18_4[7] , 
        \data_source_0/tag_data_buf_18[6]_net_1 , 
        \data_source_0/tag_data_buf_19_4[1] , 
        \data_source_0/tag_data_buf_19[0]_net_1 , 
        \data_source_0/tag_data_buf_19_4[2] , 
        \data_source_0/tag_data_buf_19[1]_net_1 , 
        \data_source_0/tag_data_buf_19_4[3] , 
        \data_source_0/tag_data_buf_19[2]_net_1 , 
        \data_source_0/tag_data_buf_19_4[4] , 
        \data_source_0/tag_data_buf_19[3]_net_1 , 
        \data_source_0/tag_data_buf_19_4[5] , 
        \data_source_0/tag_data_buf_19[4]_net_1 , 
        \data_source_0/tag_data_buf_19_4[6] , 
        \data_source_0/tag_data_buf_19[5]_net_1 , 
        \data_source_0/tag_data_buf_19_4[7] , 
        \data_source_0/tag_data_buf_19[6]_net_1 , 
        \data_source_0/tag_data_buf_20_4[1] , 
        \data_source_0/tag_data_buf_20[0]_net_1 , 
        \data_source_0/tag_data_buf_20_4[2] , 
        \data_source_0/tag_data_buf_20[1]_net_1 , 
        \data_source_0/tag_data_buf_20_4[3] , 
        \data_source_0/tag_data_buf_20[2]_net_1 , 
        \data_source_0/tag_data_buf_20_4[4] , 
        \data_source_0/tag_data_buf_20[3]_net_1 , 
        \data_source_0/tag_data_buf_20_4[5] , 
        \data_source_0/tag_data_buf_20[4]_net_1 , 
        \data_source_0/tag_data_buf_20_4[6] , 
        \data_source_0/tag_data_buf_20[5]_net_1 , 
        \data_source_0/tag_data_buf_20_4[7] , 
        \data_source_0/tag_data_buf_20[6]_net_1 , 
        \data_source_0/output_data_23[1] , 
        \data_source_0/tag_data_buf_2[7]_net_1 , 
        \data_source_0/output_data_23[3] , 
        \data_source_0/tag_data_buf_4[7]_net_1 , 
        \data_source_0/output_data_23[5] , 
        \data_source_0/tag_data_buf_6[7]_net_1 , 
        \data_source_0/output_data_23[7] , 
        \data_source_0/tag_data_buf_8[7]_net_1 , 
        \data_source_0/output_data_23[9] , 
        \data_source_0/tag_data_buf_10[7]_net_1 , 
        \data_source_0/output_data_23[11] , 
        \data_source_0/tag_data_buf_12[7]_net_1 , 
        \data_source_0/output_data_23[13] , 
        \data_source_0/tag_data_buf_14[7]_net_1 , 
        \data_source_0/output_data_23[15] , 
        \data_source_0/tag_data_buf_16[7]_net_1 , 
        \data_source_0/output_data_23[17] , 
        \data_source_0/tag_data_buf_18[7]_net_1 , 
        \data_source_0/output_data_23[19] , 
        \data_source_0/tag_data_buf_20[7]_net_1 , 
        \data_source_0/counter_n0 , \data_source_0/output_data_23[2] , 
        \data_source_0/tag_data_buf_3[7]_net_1 , 
        \data_source_0/tag_data_buf_3_4[0] , 
        \data_source_0/output_data_23[14] , 
        \data_source_0/tag_data_buf_15[7]_net_1 , 
        \data_source_0/output_data_23[6] , 
        \data_source_0/tag_data_buf_7[7]_net_1 , 
        \data_source_0/tag_data_buf_15_4[0] , 
        \data_source_0/tag_data_buf_7_4[0] , 
        \data_source_0/output_data_23[0] , 
        \data_source_0/tag_data_buf_1[7]_net_1 , 
        \data_source_0/tag_data_buf_1_4[0] , 
        \data_source_0/output_data_23[18] , 
        \data_source_0/tag_data_buf_19[7]_net_1 , 
        \data_source_0/tag_data_buf_19_4[0] , 
        \data_source_0/output_data_23[10] , 
        \data_source_0/tag_data_buf_11[7]_net_1 , 
        \data_source_0/tag_data_buf_11_4[0] , 
        \data_source_0/output_data_23[16] , 
        \data_source_0/tag_data_buf_17[7]_net_1 , 
        \data_source_0/tag_data_buf_17_4[0] , 
        \data_source_0/output_data_23[12] , 
        \data_source_0/tag_data_buf_13[7]_net_1 , 
        \data_source_0/output_data_23[4] , 
        \data_source_0/tag_data_buf_5[7]_net_1 , 
        \data_source_0/tag_data_buf_13_4[0] , 
        \data_source_0/tag_data_buf_5_4[0] , \data_source_0/N_1158 , 
        \data_source_0/N_780 , \data_source_0/N_761 , 
        \data_source_0/N_1216 , \data_source_0/N_1228 , 
        \data_source_0/N_1147 , \data_source_0/N_1150 , 
        \data_source_0/N_1221 , \data_source_0/N_758 , 
        \data_source_0/N_755 , \data_source_0/N_1020_1 , 
        \data_source_0/I_4 , \data_source_0/I_7 , \data_source_0/I_14 , 
        \data_source_0/I_17 , \data_source_0/I_23 , 
        \data_source_0/DWACT_FINC_E[2] , 
        \data_source_0/DWACT_FINC_E[3] , \data_source_0/N_3 , 
        \data_source_0/N_4 , \data_source_0/N_5 , 
        \data_source_0/DWACT_FINC_E[1] , \data_source_0/N_6 , 
        \data_source_0/N_8 , 
        \switching_circuit_0/un130_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un120_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un110_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un100_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un60_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un133_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un123_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un103_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un63_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un190_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un180_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un140_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un90_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un80_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un70_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un50_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un40_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un1_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un193_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un183_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un143_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un4_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un170_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un160_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un150_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un30_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un20_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un10_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un173_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un163_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un153_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un33_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un23_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un13_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un113_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un93_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un83_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un73_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un53_out_signal_switch_0_net_1 , 
        \switching_circuit_0/un43_out_signal_switch_0_net_1 , GND, VCC, 
        \main_clock_0/clock_out_i , \main_clock_0/counter[1]_net_1 , 
        \main_clock_0/counter[0]_net_1 , 
        \main_clock_0/counter[3]_net_1 , 
        \main_clock_0/DWACT_FINC_E[0] , \main_clock_0/counter14_4 , 
        \main_clock_0/counter14_2 , \main_clock_0/counter[2]_net_1 , 
        \main_clock_0/counter[5]_net_1 , \main_clock_0/counter14_3 , 
        \main_clock_0/counter[6]_net_1 , 
        \main_clock_0/counter[7]_net_1 , 
        \main_clock_0/counter[4]_net_1 , 
        \main_clock_0/clock_out_RNO_net_1 , 
        \main_clock_0/counter_3[0] , \main_clock_0/I_5_0 , 
        \main_clock_0/I_7_0 , \main_clock_0/I_9_0 , 
        \main_clock_0/I_12_0 , \main_clock_0/I_14_0 , 
        \main_clock_0/I_17_0 , \main_clock_0/I_20_0 , 
        \main_clock_0/N_2 , \main_clock_0/DWACT_FINC_E[2] , 
        \main_clock_0/N_3 , \main_clock_0/DWACT_FINC_E[1] , 
        \main_clock_0/N_4 , \main_clock_0/N_6 , 
        \output_signal_pad[1]/U0/NET1 , \output_signal_pad[1]/U0/NET2 , 
        \output_signal_pad[8]/U0/NET1 , \output_signal_pad[8]/U0/NET2 , 
        \output_signal_pad[13]/U0/NET1 , 
        \output_signal_pad[13]/U0/NET2 , 
        \output_signal_pad[3]/U0/NET1 , \output_signal_pad[3]/U0/NET2 , 
        \output_signal_pad[17]/U0/NET1 , 
        \output_signal_pad[17]/U0/NET2 , 
        \output_signal_pad[4]/U0/NET1 , \output_signal_pad[4]/U0/NET2 , 
        \output_signal_pad[12]/U0/NET1 , 
        \output_signal_pad[12]/U0/NET2 , 
        \output_signal_pad[19]/U0/NET1 , 
        \output_signal_pad[19]/U0/NET2 , 
        \mac_control_signal_pad/U0/NET1 , 
        \output_signal_pad[18]/U0/NET1 , 
        \output_signal_pad[18]/U0/NET2 , 
        \output_signal_pad[5]/U0/NET1 , \output_signal_pad[5]/U0/NET2 , 
        \output_signal_pad[6]/U0/NET1 , \output_signal_pad[6]/U0/NET2 , 
        \output_signal_pad[14]/U0/NET1 , 
        \output_signal_pad[14]/U0/NET2 , 
        \output_signal_pad[2]/U0/NET1 , \output_signal_pad[2]/U0/NET2 , 
        \trigger_signal_pad/U0/NET1 , \output_signal_pad[15]/U0/NET1 , 
        \output_signal_pad[15]/U0/NET2 , 
        \output_signal_pad[16]/U0/NET1 , 
        \output_signal_pad[16]/U0/NET2 , 
        \output_signal_pad[9]/U0/NET1 , \output_signal_pad[9]/U0/NET2 , 
        \output_signal_pad[10]/U0/NET1 , 
        \output_signal_pad[10]/U0/NET2 , \reset_pad/U0/NET1 , 
        \signal_into_switch_pad/U0/NET1 , 
        \signal_into_switch_pad/U0/NET2 , \clock_pad/U0/NET1 , 
        \output_signal_pad[7]/U0/NET1 , \output_signal_pad[7]/U0/NET2 , 
        \output_signal_pad[0]/U0/NET1 , \output_signal_pad[0]/U0/NET2 , 
        \output_signal_pad[11]/U0/NET1 , 
        \output_signal_pad[11]/U0/NET2 , AFLSDF_VCC, AFLSDF_GND;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign AFLSDF_GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign AFLSDF_VCC = VCC_power_net1;
    
    NOR2B \modulator_0/clock_counter_RNI41VU[11]  (.A(
        \modulator_0/clock_counter_c10 ), .B(\modulator_0/un6lto11 ), 
        .Y(\modulator_0/clock_counter_c11 ));
    DFN1E1C0 \modulator_0/clock_counter[14]  (.D(
        \modulator_0/clock_counter_n14 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/clock_counter[14]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_2_RNO[6]  (.A(
        \data_source_0/tag_data_buf_2[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_2_4[6] ));
    DFN1E1P0 \data_source_0/tag_data_buf_15[2]  (.D(
        \data_source_0/tag_data_buf_15_4[2] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_15[2]_net_1 ));
    NOR2B \data_source_0/data_index_RNID81C1[6]  (.A(
        \data_source_0/N_1211 ), .B(\data_source_0/N_1163 ), .Y(
        \data_source_0/N_860 ));
    DFN1E1C0 \data_source_0/tag_data_buf_15[4]  (.D(
        \data_source_0/tag_data_buf_15_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_15[4]_net_1 ));
    IOPAD_TRI \output_signal_pad[15]/U0/U0  (.D(
        \output_signal_pad[15]/U0/NET1 ), .E(
        \output_signal_pad[15]/U0/NET2 ), .PAD(output_signal[15]));
    OR3 \data_source_0/tag_control_sig_RNO_10[15]  (.A(
        \data_source_0/N_1056 ), .B(\data_source_0/N_1061 ), .C(
        \data_source_0/tag_control_sig_2_0_6[15] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[15] ));
    OR2A \data_source_0/tag_data_buf_5_RNO[0]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_5[7]_net_1 ), .Y(
        \data_source_0/tag_data_buf_5_4[0] ));
    NOR2B \data_source_0/tag_data_buf_4_RNO[4]  (.A(
        \data_source_0/tag_data_buf_4[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_4_4[4] ));
    MX2 \switching_circuit_0/un113_out_signal_switch_0_RNISVV51  (.A(
        \switching_circuit_0/un110_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un113_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[11] ));
    OR3 \data_source_0/tag_control_sig_RNO_2[18]  (.A(
        \data_source_0/tag_control_sig_2_0_8[18] ), .B(
        \data_source_0/tag_control_sig_2_0_7[18] ), .C(
        \data_source_0/tag_control_sig_2_0_11[18] ), .Y(
        \data_source_0/tag_control_sig_2_0_14[18] ));
    NOR2B \data_source_0/tag_data_buf_5_RNO[6]  (.A(
        \data_source_0/tag_data_buf_5[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_5_4[6] ));
    DFN1E1C0 \data_source_0/tag_data_buf_16[7]  (.D(
        \data_source_0/tag_data_buf_16_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_16[7]_net_1 ));
    OR2 \modulator_0/clock_counter_RNITDG2[7]  (.A(
        \modulator_0/clock_counter[8]_net_1 ), .B(
        \modulator_0/clock_counter[7]_net_1 ), .Y(
        \modulator_0/un6lto8 ));
    NOR2B \data_source_0/tag_control_sig_RNO_14[1]  (.A(
        \data_source_0/N_1176 ), .B(\data_source_0/N_1149 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_10_0[1] ));
    NOR3C \data_source_0/tag_control_sig_RNO_17[17]  (.A(
        \data_source_0/N_1156 ), .B(\data_source_0/N_1155 ), .C(
        \data_source_0/N_1161 ), .Y(\data_source_0/N_1100 ));
    NOR2A \data_source_0/data_index_RNI3LP8_0[1]  (.A(
        \data_source_0/data_index[1]_net_1 ), .B(
        \data_source_0/data_index[2]_net_1 ), .Y(
        \data_source_0/N_1136 ));
    IOPAD_TRI \output_signal_pad[0]/U0/U0  (.D(
        \output_signal_pad[0]/U0/NET1 ), .E(
        \output_signal_pad[0]/U0/NET2 ), .PAD(output_signal[0]));
    NOR2B \data_source_0/tag_data_buf_17_RNO[3]  (.A(
        \data_source_0/tag_data_buf_17[2]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_17_4[3] ));
    NOR2B \data_source_0/data_index_RNICN6D_2[9]  (.A(
        \data_source_0/N_1138 ), .B(
        \data_source_0/data_index[9]_net_1 ), .Y(
        \data_source_0/N_1182 ));
    DFN1E1C0 \modulator_0/clock_counter[0]  (.D(\modulator_0/N_121 ), 
        .CLK(main_clock_0_clock_out), .CLR(reset_c), .E(
        \modulator_0/clock_countere ), .Q(
        \modulator_0/clock_counter[0]_net_1 ));
    NOR3B \data_source_0/tag_control_sig_RNO_9[7]  (.A(
        \data_source_0/data_index[2]_net_1 ), .B(
        \data_source_0/tag_control_sig_2_0_a20_3_0[7] ), .C(
        \data_source_0/data_index[5]_net_1 ), .Y(\data_source_0/N_931 )
        );
    NOR3C \data_source_0/counter_RNO_1[5]  (.A(
        \data_source_0/counter[8]_net_1 ), .B(
        \data_source_0/counter[9]_net_1 ), .C(\data_source_0/N_87 ), 
        .Y(\data_source_0/N_73 ));
    NOR2A \data_source_0/data_index_RNIFQ6D_0[6]  (.A(
        \data_source_0/N_1134 ), .B(
        \data_source_0/data_index[6]_net_1 ), .Y(
        \data_source_0/N_1147 ));
    NOR2B \switching_circuit_0/un150_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[15] ), .B(
        main_clock_0_clock_out), .Y(
        \switching_circuit_0/un150_out_signal_switch_0_net_1 ));
    OR2A \data_source_0/counter_RNI9PI33[13]  (.A(
        \data_source_0/counter[13]_net_1 ), .B(\data_source_0/N_42 ), 
        .Y(\data_source_0/N_43 ));
    DFN1E1C0 \data_source_0/output_data[7]  (.D(
        \data_source_0/output_data_23[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[7] ));
    NOR2B \data_source_0/data_index_RNIIF0M_5[6]  (.A(
        \data_source_0/N_1158 ), .B(\data_source_0/N_1136 ), .Y(
        \data_source_0/N_1225 ));
    IOPAD_TRI \signal_into_switch_pad/U0/U0  (.D(
        \signal_into_switch_pad/U0/NET1 ), .E(
        \signal_into_switch_pad/U0/NET2 ), .PAD(signal_into_switch));
    NOR2B \data_source_0/tag_data_buf_7_RNO[7]  (.A(
        \data_source_0/tag_data_buf_7[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_7_4[7] ));
    DFN1E1P0 \data_source_0/tag_data_buf_14[1]  (.D(
        \data_source_0/tag_data_buf_14_4[1] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_14[1]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_10[13]  (.A(
        \data_source_0/N_1235 ), .B(\data_source_0/N_1198 ), .C(
        \data_source_0/N_1023 ), .Y(
        \data_source_0/tag_control_sig_2_0_6[13] ));
    DFN1E1P0 \data_source_0/tag_data_buf_20[4]  (.D(
        \data_source_0/tag_data_buf_20_4[4] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_20[4]_net_1 ));
    NOR2A \data_source_0/data_index_RNITJDQ[6]  (.A(
        \data_source_0/N_1162 ), .B(\data_source_0/N_701_i ), .Y(
        \data_source_0/N_919_1 ));
    OR2A \data_source_0/tag_data_buf_3_RNO[1]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_3[0]_net_1 ), .Y(
        \data_source_0/tag_data_buf_3_4[1] ));
    IOTRI_OB_EB \output_signal_pad[18]/U0/U1  (.D(
        \output_signal_c[18] ), .E(VCC), .DOUT(
        \output_signal_pad[18]/U0/NET1 ), .EOUT(
        \output_signal_pad[18]/U0/NET2 ));
    AO1 \data_source_0/tag_control_sig_RNO_4[14]  (.A(
        \data_source_0/N_729 ), .B(\data_source_0/N_1215 ), .C(
        \data_source_0/N_1038 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[14] ));
    NOR2B \data_source_0/tag_data_buf_5_RNO[4]  (.A(
        \data_source_0/tag_data_buf_5[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_5_4[4] ));
    DFN1E1 \data_source_0/tag_control_sig[1]  (.D(
        \data_source_0/tag_control_sig_2[1] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[1] ));
    AO1 \data_source_0/tag_control_sig_RNO_5[3]  (.A(
        \data_source_0/N_1200 ), .B(\data_source_0/N_1162 ), .C(
        \data_source_0/N_877 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[3] ));
    OR3 \data_source_0/tag_control_sig_RNO[1]  (.A(
        \data_source_0/tag_control_sig_2_0_12[1] ), .B(
        \data_source_0/tag_control_sig_2_0_11[1] ), .C(
        \data_source_0/tag_control_sig_2_0_16[1] ), .Y(
        \data_source_0/tag_control_sig_2[1] ));
    NOR2B \data_source_0/data_index_RNI9K6D[6]  (.A(
        \data_source_0/N_1136 ), .B(
        \data_source_0/data_index[6]_net_1 ), .Y(
        \data_source_0/N_1148 ));
    DFN1C0 \data_source_0/counter[9]  (.D(\data_source_0/N_10 ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .Q(
        \data_source_0/counter[9]_net_1 ));
    IOTRI_OB_EB \output_signal_pad[10]/U0/U1  (.D(
        \output_signal_c[10] ), .E(VCC), .DOUT(
        \output_signal_pad[10]/U0/NET1 ), .EOUT(
        \output_signal_pad[10]/U0/NET2 ));
    IOTRI_OB_EB \output_signal_pad[13]/U0/U1  (.D(
        \output_signal_c[13] ), .E(VCC), .DOUT(
        \output_signal_pad[13]/U0/NET1 ), .EOUT(
        \output_signal_pad[13]/U0/NET2 ));
    NOR2B \data_source_0/tag_control_sig_RNO_14[12]  (.A(
        \data_source_0/N_1140 ), .B(
        \data_source_0/data_index[1]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_2_1[12] ));
    XA1 \modulator_0/clock_counter_RNO[3]  (.A(
        \modulator_0/clock_counter_c2 ), .B(
        \modulator_0/clock_counter[3]_net_1 ), .C(AND2_0_Y), .Y(
        \modulator_0/clock_counter_n3 ));
    AO1 \data_source_0/tag_control_sig_RNO_14[3]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_9_0[3] ), .B(
        \data_source_0/N_1240 ), .C(\data_source_0/N_870 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[3] ));
    AND3 \main_clock_0/un5_counter_1_I_19  (.A(
        \main_clock_0/DWACT_FINC_E[0] ), .B(
        \main_clock_0/DWACT_FINC_E[2] ), .C(
        \main_clock_0/counter[6]_net_1 ), .Y(\main_clock_0/N_2 ));
    NOR2B \data_source_0/tag_data_buf_12_RNO[5]  (.A(
        \data_source_0/tag_data_buf_12[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_12_4[5] ));
    OR3 \data_source_0/tag_control_sig_RNO_0[3]  (.A(
        \data_source_0/N_867 ), .B(\data_source_0/N_876 ), .C(
        \data_source_0/tag_control_sig_2_0_3[3] ), .Y(
        \data_source_0/tag_control_sig_2_0_10[3] ));
    AND2 \data_source_0/tag_control_sig_2_0_a20_4[14]  (.A(
        \data_source_0/N_1159 ), .B(\data_source_0/N_1211 ), .Y(
        \data_source_0/N_1042 ));
    OA1 \data_source_0/tag_control_sig_RNO_6[1]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_9_0[1] ), .B(
        \data_source_0/tag_control_sig_2_0_a20_10_0[1] ), .C(
        \data_source_0/N_1156 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[1] ));
    NOR3C \data_source_0/tag_control_sig_RNO_20[3]  (.A(
        \data_source_0/N_1133 ), .B(\data_source_0/N_1151 ), .C(
        \data_source_0/N_1159 ), .Y(\data_source_0/N_870 ));
    DFN1E1C0 \data_source_0/tag_data_buf_5[1]  (.D(
        \data_source_0/tag_data_buf_5_4[1] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_5[1]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_4_RNIS3VE[7]  (.A(
        \data_source_0/tag_data_buf_4[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[3] ));
    MX2 \switching_circuit_0/out_signal_switch_1[1]  (.A(
        \switching_circuit_0/un10_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un13_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[1] ));
    OR3 \data_source_0/tag_control_sig_RNO_10[6]  (.A(
        \data_source_0/N_921 ), .B(\data_source_0/N_833 ), .C(
        \data_source_0/tag_control_sig_2_0_6[6] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[6] ));
    XA1A \switching_circuit_0/un133_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[13] ), 
        .C(\data_source_0_tag_control_sig[13] ), .Y(
        \switching_circuit_0/un133_out_signal_switch_0_net_1 ));
    NOR2B \data_source_0/tag_data_buf_8_RNO[7]  (.A(
        \data_source_0/tag_data_buf_8[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_8_4[7] ));
    XA1A \switching_circuit_0/un83_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[7] ), 
        .C(\data_source_0_tag_control_sig[8] ), .Y(
        \switching_circuit_0/un83_out_signal_switch_0_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_0[6]  (.A(
        \data_source_0/N_856 ), .B(\data_source_0/N_920 ), .C(
        \data_source_0/tag_control_sig_2_0_5[6] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[6] ));
    XA1A \data_source_0/counter_RNO[13]  (.A(\data_source_0/N_42 ), .B(
        \data_source_0/counter[13]_net_1 ), .C(
        modulator_0_output_signal), .Y(\data_source_0/counter_n13 ));
    AX1C \modulator_0/counter_RNO_0[2]  (.A(
        \modulator_0/counter[1]_net_1 ), .B(
        \modulator_0/counter[0]_net_1 ), .C(
        \modulator_0/counter[2]_net_1 ), .Y(
        \modulator_0/counter_n2_tz ));
    NOR2B \data_source_0/tag_data_buf_19_RNO[2]  (.A(
        \data_source_0/tag_data_buf_19[1]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_19_4[2] ));
    NOR2B \data_source_0/data_index_RNIIMJH_1[7]  (.A(
        \data_source_0/N_1145 ), .B(\data_source_0/N_1142 ), .Y(
        \data_source_0/N_1184 ));
    OR3 \data_source_0/tag_control_sig_RNO_4[7]  (.A(
        \data_source_0/N_939 ), .B(\data_source_0/N_927 ), .C(
        \data_source_0/tag_control_sig_2_0_4[7] ), .Y(
        \data_source_0/tag_control_sig_2_0_9[7] ));
    NOR2B \data_source_0/tag_control_sig_RNO_12[6]  (.A(
        \data_source_0/N_919_1 ), .B(\data_source_0/N_1230 ), .Y(
        \data_source_0/N_919 ));
    NOR3C \data_source_0/tag_control_sig_RNO_12[2]  (.A(
        \data_source_0/N_1133 ), .B(\data_source_0/N_1151 ), .C(
        \data_source_0/N_758 ), .Y(\data_source_0/N_849 ));
    OR2A \data_source_0/tag_data_buf_1_RNO[0]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_1[7]_net_1 ), .Y(
        \data_source_0/tag_data_buf_1_4[0] ));
    NOR2B \data_source_0/data_index_RNID81C1[4]  (.A(
        \data_source_0/N_1205 ), .B(\data_source_0/N_1163 ), .Y(
        \data_source_0/N_817 ));
    NOR2B \data_source_0/output_data_RNO[18]  (.A(
        \data_source_0/tag_data_buf_19[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[18] ));
    NOR2 \data_source_0/data_index_RNI3LP8_2[1]  (.A(
        \data_source_0/data_index[1]_net_1 ), .B(
        \data_source_0/data_index[2]_net_1 ), .Y(
        \data_source_0/N_1149 ));
    NOR3A \data_source_0/counter_RNO[5]  (.A(modulator_0_output_signal)
        , .B(\data_source_0/N_53_i ), .C(\data_source_0/N_73 ), .Y(
        \data_source_0/N_18 ));
    DFN1C0 \modulator_0/counter[2]  (.D(\modulator_0/counter_n2 ), 
        .CLK(main_clock_0_clock_out), .CLR(reset_c), .Q(
        \modulator_0/counter[2]_net_1 ));
    NOR2B \data_source_0/data_index_RNIIF0M_5[2]  (.A(
        \data_source_0/N_1155 ), .B(\data_source_0/N_1134 ), .Y(
        \data_source_0/N_1217 ));
    OR3 \data_source_0/tag_control_sig_RNO[2]  (.A(
        \data_source_0/tag_control_sig_2_0_12[2] ), .B(
        \data_source_0/tag_control_sig_2_0_11[2] ), .C(
        \data_source_0/tag_control_sig_2_0_13[2] ), .Y(
        \data_source_0/tag_control_sig_2[2] ));
    IOTRI_OB_EB \output_signal_pad[8]/U0/U1  (.D(\output_signal_c[8] ), 
        .E(VCC), .DOUT(\output_signal_pad[8]/U0/NET1 ), .EOUT(
        \output_signal_pad[8]/U0/NET2 ));
    NOR2A \data_source_0/data_index_RNIJNJH_0[7]  (.A(
        \data_source_0/N_1175 ), .B(
        \data_source_0/data_index[7]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_6_0[7] ));
    NOR3C \data_source_0/tag_control_sig_RNO_18[14]  (.A(
        \data_source_0/N_1174 ), .B(\data_source_0/N_1135 ), .C(
        \data_source_0/N_1040_1 ), .Y(\data_source_0/N_1040 ));
    NOR2B \data_source_0/tag_control_sig_RNO_6[15]  (.A(
        \data_source_0/N_1188 ), .B(\data_source_0/N_1178 ), .Y(
        \data_source_0/N_1064 ));
    NOR2B \data_source_0/tag_data_buf_8_RNO[1]  (.A(
        \data_source_0/tag_data_buf_8[0]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_8_4[1] ));
    DFN1E1C0 \data_source_0/tag_data_buf_1[1]  (.D(
        \data_source_0/tag_data_buf_1_4[1] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_1[1]_net_1 ));
    OR2 \data_source_0/tag_control_sig_RNO_19[4]  (.A(
        \data_source_0/N_1186 ), .B(\data_source_0/N_1162 ), .Y(
        \data_source_0/N_534_tz ));
    OR3 \data_source_0/tag_control_sig_RNO[5]  (.A(
        \data_source_0/tag_control_sig_2_0_12[5] ), .B(
        \data_source_0/tag_control_sig_2_0_11[5] ), .C(
        \data_source_0/tag_control_sig_2_0_13[5] ), .Y(
        \data_source_0/tag_control_sig_2[5] ));
    NOR3C \data_source_0/tag_control_sig_RNO_12[11]  (.A(
        \data_source_0/N_1148 ), .B(
        \data_source_0/data_index_0[4]_net_1 ), .C(
        \data_source_0/N_1184 ), .Y(\data_source_0/N_995 ));
    NOR2B \data_source_0/data_index_RNIU6731[9]  (.A(
        \data_source_0/N_1211 ), .B(\data_source_0/N_1175 ), .Y(
        \data_source_0/N_921 ));
    DFN1E1P0 \data_source_0/tag_data_buf_14[3]  (.D(
        \data_source_0/tag_data_buf_14_4[3] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_14[3]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_17[6]  (.A(
        \data_source_0/N_1242 ), .B(\data_source_0/N_1187 ), .C(
        \data_source_0/N_925 ), .Y(
        \data_source_0/tag_control_sig_2_0_6[6] ));
    DFN1E1 \data_source_0/tag_control_sig[15]  (.D(
        \data_source_0/tag_control_sig_2[15] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[15] ));
    NOR2B \data_source_0/tag_data_buf_17_RNO[2]  (.A(
        \data_source_0/tag_data_buf_17[1]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_17_4[2] ));
    OR3 \data_source_0/tag_control_sig_RNO_0[14]  (.A(
        \data_source_0/tag_control_sig_2_0_1[14] ), .B(
        \data_source_0/tag_control_sig_2_0_0[14] ), .C(
        \data_source_0/tag_control_sig_2_0_8[14] ), .Y(
        \data_source_0/tag_control_sig_2_0_13[14] ));
    NOR3C \data_source_0/tag_control_sig_RNO_13[8]  (.A(
        \data_source_0/N_1156 ), .B(\data_source_0/N_1155 ), .C(
        \data_source_0/N_1141 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_10_0[8] ));
    OR3 \data_source_0/tag_control_sig_RNO_10[10]  (.A(
        \data_source_0/N_978 ), .B(\data_source_0/N_979 ), .C(
        \data_source_0/tag_control_sig_2_0_4[10] ), .Y(
        \data_source_0/tag_control_sig_2_0_9[10] ));
    NOR3C \data_source_0/tag_control_sig_RNO_13[11]  (.A(
        \data_source_0/N_1178 ), .B(\data_source_0/N_1156 ), .C(
        \data_source_0/N_1233 ), .Y(\data_source_0/N_988 ));
    DFN1E1 \data_source_0/tag_control_sig[17]  (.D(
        \data_source_0/tag_control_sig_2[17] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[17] ));
    NOR2B \data_source_0/data_index_RNIIF0M_2[2]  (.A(
        \data_source_0/N_1157 ), .B(\data_source_0/N_1156 ), .Y(
        \data_source_0/N_1216 ));
    DFN1E1C0 \data_source_0/tag_data_buf_8[6]  (.D(
        \data_source_0/tag_data_buf_8_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_8[6]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_8[1]  (.A(
        \data_source_0/N_1207 ), .B(\data_source_0/N_1182 ), .C(
        \data_source_0/N_837 ), .Y(
        \data_source_0/tag_control_sig_2_0_4[1] ));
    IOTRI_OB_EB \output_signal_pad[4]/U0/U1  (.D(\output_signal_c[4] ), 
        .E(VCC), .DOUT(\output_signal_pad[4]/U0/NET1 ), .EOUT(
        \output_signal_pad[4]/U0/NET2 ));
    DFN1E1C0 \data_source_0/tag_data_buf_16[1]  (.D(
        \data_source_0/tag_data_buf_16_4[1] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_16[1]_net_1 ));
    XOR2 \data_source_0/data_index_RNIBTP8[6]  (.A(
        \data_source_0/data_index[6]_net_1 ), .B(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/N_701_i ));
    NOR2B \data_source_0/tag_control_sig_RNO_14[0]  (.A(
        \data_source_0/N_1216 ), .B(\data_source_0/N_1162 ), .Y(
        \data_source_0/N_823 ));
    DFN1E1C0 \data_source_0/tag_data_buf_7[5]  (.D(
        \data_source_0/tag_data_buf_7_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_7[5]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_4[5]  (.D(
        \data_source_0/tag_data_buf_4_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_4[5]_net_1 ));
    IOPAD_IN \reset_pad/U0/U0  (.PAD(reset), .Y(\reset_pad/U0/NET1 ));
    NOR2B \data_source_0/tag_data_buf_1_RNO[2]  (.A(
        \data_source_0/tag_data_buf_1[1]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_1_4[2] ));
    NOR2B \data_source_0/tag_control_sig_RNO_24[1]  (.A(
        \data_source_0/N_1197 ), .B(\data_source_0/N_1181 ), .Y(
        \data_source_0/N_846 ));
    NOR2B \data_source_0/data_index_RNIIF0M_3[6]  (.A(
        \data_source_0/N_1158 ), .B(\data_source_0/N_1149 ), .Y(
        \data_source_0/N_1188 ));
    NOR2B \data_source_0/tag_data_buf_14_RNO[5]  (.A(
        \data_source_0/tag_data_buf_14[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_14_4[5] ));
    NOR3C \data_source_0/tag_control_sig_RNO_15[8]  (.A(
        \data_source_0/N_1140 ), .B(\data_source_0/N_1154 ), .C(
        \data_source_0/N_1177 ), .Y(\data_source_0/N_952 ));
    XA1A \switching_circuit_0/un63_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[6] ), 
        .C(\data_source_0_tag_control_sig[6] ), .Y(
        \switching_circuit_0/un63_out_signal_switch_0_net_1 ));
    NOR2B \data_source_0/output_data_RNO[6]  (.A(
        \data_source_0/tag_data_buf_7[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[6] ));
    NOR2B \data_source_0/data_index_RNI7PP8_0[5]  (.A(
        \data_source_0/data_index[2]_net_1 ), .B(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/N_1228 ));
    DFN1E1C0 \data_source_0/tag_data_buf_19[5]  (.D(
        \data_source_0/tag_data_buf_19_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_19[5]_net_1 ));
    XOR2 \main_clock_0/un5_counter_1_I_9  (.A(\main_clock_0/N_6 ), .B(
        \main_clock_0/counter[3]_net_1 ), .Y(\main_clock_0/I_9_0 ));
    DFN1E1C0 \data_source_0/tag_data_buf_6[5]  (.D(
        \data_source_0/tag_data_buf_6_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_6[5]_net_1 ));
    NOR2B \data_source_0/data_index_RNIIF0M_0[4]  (.A(
        \data_source_0/N_1154 ), .B(\data_source_0/N_1134 ), .Y(
        \data_source_0/N_1205 ));
    NOR3 \data_source_0/counter_RNIRCTA[15]  (.A(
        \data_source_0/counter[5]_net_1 ), .B(
        \data_source_0/counter[15]_net_1 ), .C(
        \data_source_0/counter[12]_net_1 ), .Y(
        \data_source_0/counter_n9_i_a2_4 ));
    AO1 \data_source_0/tag_control_sig_RNO_7[4]  (.A(
        \data_source_0/N_1183 ), .B(\data_source_0/N_1180 ), .C(
        \data_source_0/N_888 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[4] ));
    OR2A \data_source_0/tag_data_buf_12_RNO[3]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_12[2]_net_1 ), .Y(
        \data_source_0/tag_data_buf_12_4[3] ));
    NOR2B \data_source_0/tag_control_sig_RNO_21[17]  (.A(
        \data_source_0/N_1123_1 ), .B(\data_source_0/N_1177 ), .Y(
        \data_source_0/N_1096 ));
    NOR3B \data_source_0/tag_control_sig_RNO_12[0]  (.A(
        \data_source_0/N_1185 ), .B(\data_source_0/N_813_1 ), .C(
        \data_source_0/N_707_i ), .Y(\data_source_0/N_813 ));
    DFN1C0 \data_source_0/data_index[7]  (.D(
        \data_source_0/data_index_3[7] ), .CLK(
        modulator_0_output_signal), .CLR(reset_c), .Q(
        \data_source_0/data_index[7]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_9[3]  (.A(
        \data_source_0/N_879 ), .B(\data_source_0/N_875 ), .C(
        \data_source_0/tag_control_sig_2_0_5[3] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[3] ));
    AO1 \data_source_0/tag_control_sig_RNO_7[10]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_3_1[10] ), .B(
        \data_source_0/tag_control_sig_2_0_a20_3_0[10] ), .C(
        \data_source_0/N_981 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[10] ));
    AO1 \data_source_0/tag_control_sig_RNO_22[18]  (.A(
        \data_source_0/N_1189 ), .B(\data_source_0/N_1159 ), .C(
        \data_source_0/N_1103 ), .Y(
        \data_source_0/tag_control_sig_2_0_6[18] ));
    NOR2B \data_source_0/data_index_RNIIF0M_1[5]  (.A(
        \data_source_0/N_1150 ), .B(\data_source_0/N_1149 ), .Y(
        \data_source_0/N_1183 ));
    DFN1E1C0 \modulator_0/clock_counter[2]  (.D(
        \modulator_0/clock_counter_n2 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/clock_counter[2]_net_1 ));
    NOR2B \switching_circuit_0/un190_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[19] ), .B(
        main_clock_0_clock_out), .Y(
        \switching_circuit_0/un190_out_signal_switch_0_net_1 ));
    NOR3C \modulator_0/counter_RNO_0[5]  (.A(
        \modulator_0/counter[3]_net_1 ), .B(\modulator_0/counter_c2 ), 
        .C(\modulator_0/counter[4]_net_1 ), .Y(
        \modulator_0/counter_45_0 ));
    DFN1C0 \main_clock_0/counter[1]  (.D(\main_clock_0/I_5_0 ), .CLK(
        GLA), .CLR(reset_c), .Q(\main_clock_0/counter[1]_net_1 ));
    NOR2B \data_source_0/data_index_RNID81C1[5]  (.A(
        \data_source_0/N_1204 ), .B(\data_source_0/N_1176 ), .Y(
        \data_source_0/N_903 ));
    NOR2B \data_source_0/tag_control_sig_RNO_16[11]  (.A(
        \data_source_0/N_1206 ), .B(\data_source_0/N_1159 ), .Y(
        \data_source_0/N_993 ));
    NOR2A \data_source_0/tag_control_sig_RNO_23[18]  (.A(
        \data_source_0/N_1152 ), .B(
        \data_source_0/data_index[4]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_4_1[18] ));
    OR3 \data_source_0/tag_control_sig_RNO_10[2]  (.A(
        \data_source_0/N_1220 ), .B(\data_source_0/N_1219 ), .C(
        \data_source_0/N_764 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[2] ));
    OR2 \data_source_0/data_index_RNI4V0C1_0[2]  (.A(
        \data_source_0/N_1210 ), .B(\data_source_0/N_1197 ), .Y(
        \data_source_0/N_757 ));
    NOR2B \data_source_0/tag_data_buf_11_RNO[5]  (.A(
        \data_source_0/tag_data_buf_11[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_11_4[5] ));
    NOR2B \modulator_0/clock_counter_RNIFVF2[1]  (.A(
        \modulator_0/clock_counter[1]_net_1 ), .B(
        \modulator_0/clock_counter[0]_net_1 ), .Y(
        \modulator_0/clock_counter_c1 ));
    AO1 \data_source_0/tag_control_sig_RNO_9[14]  (.A(
        \data_source_0/N_802 ), .B(\data_source_0/N_1189 ), .C(
        \data_source_0/N_1052 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[14] ));
    OR3 \data_source_0/tag_control_sig_RNO_2[8]  (.A(
        \data_source_0/tag_control_sig_2_0_5[8] ), .B(
        \data_source_0/tag_control_sig_2_0_4[8] ), .C(
        \data_source_0/tag_control_sig_2_0_11[8] ), .Y(
        \data_source_0/tag_control_sig_2_0_13[8] ));
    XA1 \modulator_0/clock_counter_RNO[7]  (.A(
        \modulator_0/clock_counter_c6 ), .B(
        \modulator_0/clock_counter[7]_net_1 ), .C(AND2_0_Y), .Y(
        \modulator_0/clock_counter_n7 ));
    DFN1E1C0 \data_source_0/tag_data_buf_3[7]  (.D(
        \data_source_0/tag_data_buf_3_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_3[7]_net_1 ));
    AO1 \data_source_0/tag_control_sig_2_0_7[11]  (.A(
        \data_source_0/N_1159 ), .B(\data_source_0/N_1196 ), .C(
        \data_source_0/N_994 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[11]_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_16[1]  (.A(
        \data_source_0/N_1133 ), .B(\data_source_0/N_1151 ), .C(
        \data_source_0/N_1177 ), .Y(\data_source_0/N_834 ));
    DFN1E1C0 \data_source_0/tag_data_buf_8[0]  (.D(
        \data_source_0/output_data_23[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_8[0]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_8[3]  (.A(
        \data_source_0/N_1202 ), .B(\data_source_0/N_1163 ), .C(
        \data_source_0/N_869 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[3] ));
    NOR2B \data_source_0/data_index_RNIIMJH_0[0]  (.A(
        \data_source_0/N_1145 ), .B(\data_source_0/N_1138 ), .Y(
        \data_source_0/N_1174 ));
    NOR2B \modulator_0/clock_counter_RNI6GO8[6]  (.A(
        \modulator_0/clock_counter_c5 ), .B(\modulator_0/un5lto6 ), .Y(
        \modulator_0/clock_counter_c6 ));
    NOR2B \data_source_0/tag_data_buf_18_RNO[6]  (.A(
        \data_source_0/tag_data_buf_18[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_18_4[6] ));
    DFN1E1C0 \data_source_0/tag_data_buf_16[0]  (.D(
        \data_source_0/output_data_23[15] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_16[0]_net_1 ));
    DFN1E1C0 \modulator_0/clock_counter[11]  (.D(
        \modulator_0/clock_counter_n11 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/un6lto11 ));
    AO1 \data_source_0/tag_control_sig_RNO_18[18]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_4_1[18] ), .B(
        \data_source_0/tag_control_sig_2_0_a20_4_0[18] ), .C(
        \data_source_0/N_1027 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[18] ));
    NOR2B \data_source_0/tag_control_sig_RNO_20[6]  (.A(
        \data_source_0/N_1210 ), .B(\data_source_0/N_1161 ), .Y(
        \data_source_0/N_925 ));
    NOR2B \data_source_0/data_index_RNIIF0M_6[6]  (.A(
        \data_source_0/N_1158 ), .B(\data_source_0/N_1152 ), .Y(
        \data_source_0/N_1235 ));
    NOR2B \data_source_0/tag_control_sig_RNO_17[5]  (.A(
        \data_source_0/N_807 ), .B(\data_source_0/N_1188 ), .Y(
        \data_source_0/N_897 ));
    AO1 \data_source_0/tag_control_sig_RNO_5[14]  (.A(
        \data_source_0/N_1209 ), .B(\data_source_0/N_1177 ), .C(
        \data_source_0/N_1046 ), .Y(
        \data_source_0/tag_control_sig_2_0_8[14] ));
    OA1 \data_source_0/tag_control_sig_RNO_19[7]  (.A(
        \data_source_0/N_1227 ), .B(\data_source_0/N_1232 ), .C(
        \data_source_0/N_1179 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_3_0[7] ));
    DFN1E1C0 \data_source_0/tag_data_buf_4[4]  (.D(
        \data_source_0/tag_data_buf_4_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_4[4]_net_1 ));
    OR3 \modulator_0/output_signal_RNO_5  (.A(\modulator_0/un5lto15_2 )
        , .B(\modulator_0/un5lto15_1 ), .C(\modulator_0/un5lto15_3 ), 
        .Y(\modulator_0/un5lto15_6 ));
    OR2A \data_source_0/tag_data_buf_19_RNO[4]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_19[3]_net_1 ), .Y(
        \data_source_0/tag_data_buf_19_4[4] ));
    NOR3A \data_source_0/counter_RNI2O3C[13]  (.A(
        \data_source_0/counter_n9_i_a2_4 ), .B(
        \data_source_0/counter[14]_net_1 ), .C(
        \data_source_0/counter[13]_net_1 ), .Y(
        \data_source_0/counter_n9_i_a2_6 ));
    OR2A \data_source_0/tag_data_buf_16_RNO[4]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_16[3]_net_1 ), .Y(
        \data_source_0/tag_data_buf_16_4[4] ));
    OR2A \data_source_0/tag_data_buf_11_RNO[0]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_11[7]_net_1 ), .Y(
        \data_source_0/tag_data_buf_11_4[0] ));
    NOR2 \data_source_0/data_index_RNI3LP8_3[0]  (.A(
        \data_source_0/data_index[0]_net_1 ), .B(
        \data_source_0/data_index[3]_net_1 ), .Y(
        \data_source_0/N_1141 ));
    XA1 \modulator_0/clock_counter_RNO[8]  (.A(
        \modulator_0/clock_counter_c7 ), .B(
        \modulator_0/clock_counter[8]_net_1 ), .C(AND2_0_Y), .Y(
        \modulator_0/clock_counter_n8 ));
    DFN1E1 \data_source_0/tag_control_sig[19]  (.D(
        \data_source_0/tag_control_sig_2[19] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[19] ));
    DFN1C0 \data_source_0/counter[5]  (.D(\data_source_0/N_18 ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .Q(
        \data_source_0/counter[5]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_8[7]  (.D(
        \data_source_0/tag_data_buf_8_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_8[7]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_26[18]  (.A(
        \data_source_0/N_755 ), .B(\data_source_0/N_1216 ), .Y(
        \data_source_0/N_1103 ));
    IOTRI_OB_EB \output_signal_pad[0]/U0/U1  (.D(\output_signal_c[0] ), 
        .E(VCC), .DOUT(\output_signal_pad[0]/U0/NET1 ), .EOUT(
        \output_signal_pad[0]/U0/NET2 ));
    DFN1E1C0 \data_source_0/tag_data_buf_8[4]  (.D(
        \data_source_0/tag_data_buf_8_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_8[4]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_2[5]  (.A(
        \data_source_0/tag_control_sig_2_0_4[5] ), .B(
        \data_source_0/tag_control_sig_2_0_3[5] ), .C(
        \data_source_0/tag_control_sig_2_0_9[5] ), .Y(
        \data_source_0/tag_control_sig_2_0_13[5] ));
    DFN1E1C0 \data_source_0/tag_data_buf_18[0]  (.D(
        \data_source_0/output_data_23[17] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_18[0]_net_1 ));
    NOR3B \data_source_0/tag_control_sig_RNO_7[17]  (.A(
        \data_source_0/N_1160 ), .B(\data_source_0/N_1230 ), .C(
        \data_source_0/N_701_i ), .Y(\data_source_0/N_1090 ));
    AO1 \data_source_0/tag_control_sig_RNO_5[1]  (.A(
        \data_source_0/N_1209 ), .B(\data_source_0/N_1198 ), .C(
        \data_source_0/N_841 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[1] ));
    NOR2B \data_source_0/tag_control_sig_RNO_11[3]  (.A(
        \data_source_0/N_1187 ), .B(\data_source_0/N_1179 ), .Y(
        \data_source_0/N_877 ));
    NOR2B \data_source_0/tag_data_buf_20_RNO[5]  (.A(
        \data_source_0/tag_data_buf_20[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_20_4[5] ));
    NOR2B \data_source_0/tag_control_sig_RNO_13[1]  (.A(
        \data_source_0/N_1162 ), .B(\data_source_0/N_1133 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_9_0[1] ));
    DFN1E1C0 \data_source_0/output_data[1]  (.D(
        \data_source_0/output_data_23[1] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[1] ));
    DFN1E1P0 \data_source_0/tag_data_buf_7[2]  (.D(
        \data_source_0/tag_data_buf_7_4[2] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_7[2]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_13[12]  (.A(
        \data_source_0/N_1201 ), .B(\data_source_0/N_1162 ), .Y(
        \data_source_0/N_1014 ));
    IOPAD_IN \trigger_signal_pad/U0/U0  (.PAD(trigger_signal), .Y(
        \trigger_signal_pad/U0/NET1 ));
    MX2 \switching_circuit_0/out_signal_switch_1[10]  (.A(
        \switching_circuit_0/un100_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un103_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[10] ));
    DFN1C0 \data_source_0/data_index[5]  (.D(\data_source_0/I_14 ), 
        .CLK(modulator_0_output_signal), .CLR(reset_c), .Q(
        \data_source_0/data_index[5]_net_1 ));
    IOPAD_TRI \output_signal_pad[14]/U0/U0  (.D(
        \output_signal_pad[14]/U0/NET1 ), .E(
        \output_signal_pad[14]/U0/NET2 ), .PAD(output_signal[14]));
    NOR3C \data_source_0/data_index_RNIJ6UA1[2]  (.A(
        \data_source_0/N_1156 ), .B(\data_source_0/N_1155 ), .C(
        \data_source_0/N_1180 ), .Y(\data_source_0/N_872 ));
    OR2A \data_source_0/tag_data_buf_20_RNO[4]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_20[3]_net_1 ), .Y(
        \data_source_0/tag_data_buf_20_4[4] ));
    PLLBA \pll_core_0/Core  (.CLKA(clock_c), .EXTFB(GND), .POWERDOWN(
        VCC), .GLA(GLA), .LOCK(), .GLB(), .YB(), .GLC(), .YC(), 
        .OADIV0(GND), .OADIV1(GND), .OADIV2(GND), .OADIV3(GND), 
        .OADIV4(GND), .OAMUX0(GND), .OAMUX1(GND), .OAMUX2(VCC), 
        .DLYGLA0(GND), .DLYGLA1(GND), .DLYGLA2(GND), .DLYGLA3(GND), 
        .DLYGLA4(GND), .OBDIV0(AFLSDF_GND), .OBDIV1(AFLSDF_GND), 
        .OBDIV2(AFLSDF_GND), .OBDIV3(AFLSDF_GND), .OBDIV4(AFLSDF_GND), 
        .OBMUX0(AFLSDF_GND), .OBMUX1(AFLSDF_GND), .OBMUX2(AFLSDF_GND), 
        .DLYYB0(AFLSDF_GND), .DLYYB1(AFLSDF_GND), .DLYYB2(AFLSDF_GND), 
        .DLYYB3(AFLSDF_GND), .DLYYB4(AFLSDF_GND), .DLYGLB0(AFLSDF_GND), 
        .DLYGLB1(AFLSDF_GND), .DLYGLB2(AFLSDF_GND), .DLYGLB3(
        AFLSDF_GND), .DLYGLB4(AFLSDF_GND), .OCDIV0(AFLSDF_GND), 
        .OCDIV1(AFLSDF_GND), .OCDIV2(AFLSDF_GND), .OCDIV3(AFLSDF_GND), 
        .OCDIV4(AFLSDF_GND), .OCMUX0(AFLSDF_GND), .OCMUX1(AFLSDF_GND), 
        .OCMUX2(AFLSDF_GND), .DLYYC0(AFLSDF_GND), .DLYYC1(AFLSDF_GND), 
        .DLYYC2(AFLSDF_GND), .DLYYC3(AFLSDF_GND), .DLYYC4(AFLSDF_GND), 
        .DLYGLC0(AFLSDF_GND), .DLYGLC1(AFLSDF_GND), .DLYGLC2(
        AFLSDF_GND), .DLYGLC3(AFLSDF_GND), .DLYGLC4(AFLSDF_GND), 
        .FINDIV0(VCC), .FINDIV1(VCC), .FINDIV2(GND), .FINDIV3(GND), 
        .FINDIV4(GND), .FINDIV5(GND), .FINDIV6(GND), .FBDIV0(VCC), 
        .FBDIV1(VCC), .FBDIV2(GND), .FBDIV3(GND), .FBDIV4(VCC), 
        .FBDIV5(GND), .FBDIV6(GND), .FBDLY0(GND), .FBDLY1(GND), 
        .FBDLY2(GND), .FBDLY3(GND), .FBDLY4(GND), .FBSEL0(VCC), 
        .FBSEL1(GND), .XDLYSEL(GND), .VCOSEL0(GND), .VCOSEL1(GND), 
        .VCOSEL2(VCC));
    NOR3B \data_source_0/data_index_0_RNI1NTK_2[7]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/N_1142 ), .C(
        \data_source_0/data_index_0[7]_net_1 ), .Y(
        \data_source_0/N_1185 ));
    NOR2B \switching_circuit_0/un10_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[1] ), .B(main_clock_0_clock_out)
        , .Y(\switching_circuit_0/un10_out_signal_switch_0_net_1 ));
    NOR2B \data_source_0/data_index_RNIIF0M_4[2]  (.A(
        \data_source_0/N_1155 ), .B(\data_source_0/N_1140 ), .Y(
        \data_source_0/N_1199 ));
    MX2 \switching_circuit_0/out_signal_switch_1[2]  (.A(
        \switching_circuit_0/un20_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un23_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[2] ));
    NOR2B \data_source_0/tag_data_buf_11_RNO[2]  (.A(
        \data_source_0/tag_data_buf_11[1]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_11_4[2] ));
    NOR2B \data_source_0/tag_data_buf_10_RNO[2]  (.A(
        \data_source_0/tag_data_buf_10[1]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_10_4[2] ));
    DFN1E1C0 \modulator_0/clock_counter[13]  (.D(
        \modulator_0/clock_counter_n13 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/clock_counter[13]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_3[3]  (.D(
        \data_source_0/tag_data_buf_3_4[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_3[3]_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_21[14]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/N_1141 ), .C(\data_source_0/N_1183 ), .Y(
        \data_source_0/N_1045 ));
    OR2 \data_source_0/tag_control_sig_RNO_22[12]  (.A(
        \data_source_0/N_1208 ), .B(\data_source_0/N_1134 ), .Y(
        \data_source_0/N_771 ));
    NOR2B \data_source_0/tag_data_buf_3_RNO[2]  (.A(
        \data_source_0/tag_data_buf_3[1]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_3_4[2] ));
    OA1 \data_source_0/data_index_RNIT5731[5]  (.A(
        \data_source_0/N_1227 ), .B(\data_source_0/N_1232 ), .C(
        \data_source_0/N_1228 ), .Y(\data_source_0/N_1244 ));
    NOR2B \data_source_0/tag_control_sig_RNO_22[15]  (.A(
        \data_source_0/N_1134 ), .B(
        \data_source_0/data_index[2]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_0_1[15] ));
    OR3 \data_source_0/tag_control_sig_RNO[9]  (.A(
        \data_source_0/tag_control_sig_2_0_13[9] ), .B(
        \data_source_0/tag_control_sig_2_0_12[9] ), .C(
        \data_source_0/tag_control_sig_2_0_14[9] ), .Y(
        \data_source_0/tag_control_sig_2[9] ));
    OR3 \data_source_0/tag_control_sig_RNO[18]  (.A(
        \data_source_0/tag_control_sig_2_0_10[18] ), .B(
        \data_source_0/tag_control_sig_2_0_9[18] ), .C(
        \data_source_0/tag_control_sig_2_0_14[18] ), .Y(
        \data_source_0/tag_control_sig_2[18] ));
    DFN1E1C0 \data_source_0/tag_data_buf_17[3]  (.D(
        \data_source_0/tag_data_buf_17_4[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_17[3]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO[6]  (.A(
        \data_source_0/tag_control_sig_2_0_11[6] ), .B(
        \data_source_0/tag_control_sig_2_0_10[6] ), .C(
        \data_source_0/tag_control_sig_2_0_15[6] ), .Y(
        \data_source_0/tag_control_sig_2[6] ));
    NOR2B \data_source_0/tag_control_sig_RNO_13[9]  (.A(
        \data_source_0/N_1190 ), .B(\data_source_0/N_1162 ), .Y(
        \data_source_0/N_964 ));
    AO1 \modulator_0/output_signal_RNO_4  (.A(\modulator_0/un5lto5 ), 
        .B(\modulator_0/un5lto6 ), .C(\modulator_0/un6lto8 ), .Y(
        \modulator_0/un5lto15_5 ));
    NOR2B \data_source_0/tag_control_sig_RNO_23[15]  (.A(
        \data_source_0/N_1187 ), .B(\data_source_0/N_1176 ), .Y(
        \data_source_0/N_1059 ));
    DFN1E1C0 \data_source_0/output_data[2]  (.D(
        \data_source_0/output_data_23[2] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[2] ));
    AND2 \data_source_0/un3_data_index_I_15  (.A(
        \data_source_0/data_index[3]_net_1 ), .B(
        \data_source_0/data_index_0[4]_net_1 ), .Y(
        \data_source_0/DWACT_FINC_E[1] ));
    DFN1C0 \data_source_0/counter[12]  (.D(\data_source_0/counter_n12 )
        , .CLK(main_clock_0_clock_out), .CLR(reset_c), .Q(
        \data_source_0/counter[12]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_17[5]  (.D(
        \data_source_0/tag_data_buf_17_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_17[5]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_13_RNO[5]  (.A(
        \data_source_0/tag_data_buf_13[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_13_4[5] ));
    NOR3B \data_source_0/data_index_0_RNI9A421[4]  (.A(
        \data_source_0/N_1159 ), .B(\data_source_0/N_1136 ), .C(
        \data_source_0/N_759 ), .Y(\data_source_0/N_904 ));
    NOR2B \data_source_0/tag_data_buf_4_RNO[6]  (.A(
        \data_source_0/tag_data_buf_4[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_4_4[6] ));
    OR2A \data_source_0/tag_data_buf_19_RNO[1]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_19[0]_net_1 ), .Y(
        \data_source_0/tag_data_buf_19_4[1] ));
    NOR2B \data_source_0/tag_data_buf_16_RNO[2]  (.A(
        \data_source_0/tag_data_buf_16[1]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_16_4[2] ));
    OA1 \data_source_0/tag_control_sig_RNO_16[12]  (.A(
        \data_source_0/N_1187 ), .B(\data_source_0/N_1201 ), .C(
        \data_source_0/N_1184 ), .Y(\data_source_0/N_1007 ));
    NOR2B \data_source_0/tag_data_buf_10_RNO[6]  (.A(
        \data_source_0/tag_data_buf_10[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_10_4[6] ));
    NOR2B \data_source_0/tag_data_buf_6_RNO[6]  (.A(
        \data_source_0/tag_data_buf_6[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_6_4[6] ));
    NOR3C \data_source_0/tag_control_sig_RNO_19[11]  (.A(
        \data_source_0/N_1142 ), .B(\data_source_0/N_1139 ), .C(
        \data_source_0/N_1188 ), .Y(\data_source_0/N_997 ));
    NOR2B \data_source_0/counter_RNO_1[8]  (.A(
        \data_source_0/counter[9]_net_1 ), .B(\data_source_0/N_87 ), 
        .Y(\data_source_0/counter_n8_i_a3_0_0 ));
    AO1 \data_source_0/tag_control_sig_RNO_5[5]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_3_0[5] ), .B(
        \data_source_0/N_901_1 ), .C(\data_source_0/N_911 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[5] ));
    NOR2B \data_source_0/tag_control_sig_RNO_17[2]  (.A(
        \data_source_0/N_1188 ), .B(\data_source_0/N_1175 ), .Y(
        \data_source_0/N_854 ));
    AO1 \data_source_0/tag_control_sig_RNO_6[19]  (.A(
        \data_source_0/N_1207 ), .B(\data_source_0/N_1177 ), .C(
        \data_source_0/tag_control_sig_RNO_12[19]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[19] ));
    AO1 \data_source_0/tag_control_sig_RNO_10[14]  (.A(
        \data_source_0/N_1195 ), .B(\data_source_0/N_1182 ), .C(
        \data_source_0/N_1050 ), .Y(
        \data_source_0/tag_control_sig_2_0_4[14] ));
    OR2A \data_source_0/tag_data_buf_12_RNO[2]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_12[1]_net_1 ), .Y(
        \data_source_0/tag_data_buf_12_4[2] ));
    AO1 \modulator_0/output_signal_RNO_6  (.A(\modulator_0/un6lto6_0 ), 
        .B(\modulator_0/un6lto4 ), .C(\modulator_0/un6lto8 ), .Y(
        \modulator_0/un6lt9 ));
    OR3 \data_source_0/tag_control_sig_RNO_1[2]  (.A(
        \data_source_0/N_863 ), .B(\data_source_0/N_862 ), .C(
        \data_source_0/tag_control_sig_2_0_6[2] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[2] ));
    DFN1E1 \data_source_0/tag_control_sig[11]  (.D(
        \data_source_0/tag_control_sig_2[11] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[11] ));
    DFN1E1C0 \data_source_0/tag_data_buf_20[7]  (.D(
        \data_source_0/tag_data_buf_20_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_20[7]_net_1 ));
    OR2 \data_source_0/tag_control_sig_RNO_12[3]  (.A(
        \data_source_0/N_1182 ), .B(\data_source_0/N_1181 ), .Y(
        \data_source_0/N_808 ));
    AO1 \data_source_0/tag_control_sig_RNO_7[18]  (.A(
        \data_source_0/N_1188 ), .B(\data_source_0/N_1180 ), .C(
        \data_source_0/N_1115 ), .Y(
        \data_source_0/tag_control_sig_2_0_2[18] ));
    NOR2B \data_source_0/tag_data_buf_5_RNO[1]  (.A(
        \data_source_0/tag_data_buf_5[0]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_5_4[1] ));
    NOR2B \data_source_0/tag_control_sig_RNO_8[7]  (.A(
        \data_source_0/N_1210 ), .B(\data_source_0/N_1160 ), .Y(
        \data_source_0/N_935 ));
    NOR2B \data_source_0/data_index_RNIIMJH_1[0]  (.A(
        \data_source_0/N_1141 ), .B(\data_source_0/N_1144 ), .Y(
        \data_source_0/N_1178 ));
    MX2 \switching_circuit_0/out_signal_switch_1[16]  (.A(
        \switching_circuit_0/un160_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un163_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[16] ));
    DFN1C0 \data_source_0/data_index[2]  (.D(\data_source_0/I_7 ), 
        .CLK(modulator_0_output_signal), .CLR(reset_c), .Q(
        \data_source_0/data_index[2]_net_1 ));
    DFN1C0 \main_clock_0/clock_out  (.D(
        \main_clock_0/clock_out_RNO_net_1 ), .CLK(GLA), .CLR(reset_c), 
        .Q(\main_clock_0/clock_out_i ));
    DFN1E1C0 \data_source_0/tag_data_buf_15[5]  (.D(
        \data_source_0/tag_data_buf_15_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_15[5]_net_1 ));
    OA1 \data_source_0/tag_control_sig_RNO_14[2]  (.A(
        \data_source_0/N_1187 ), .B(\data_source_0/N_1201 ), .C(
        \data_source_0/N_1174 ), .Y(\data_source_0/N_851 ));
    DFN1E1C0 \modulator_0/clock_counter[3]  (.D(
        \modulator_0/clock_counter_n3 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/clock_counter[3]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_6[12]  (.A(
        \data_source_0/N_1235 ), .B(\data_source_0/N_1179 ), .Y(
        \data_source_0/N_1018 ));
    NOR2A \data_source_0/data_index_RNI9RP8_0[4]  (.A(
        \data_source_0/data_index[5]_net_1 ), .B(
        \data_source_0/data_index[4]_net_1 ), .Y(
        \data_source_0/N_1156 ));
    OR3 \data_source_0/tag_control_sig_RNO_7[7]  (.A(
        \data_source_0/N_930 ), .B(\data_source_0/N_929 ), .C(
        \data_source_0/tag_control_sig_2_0_1[7] ), .Y(
        \data_source_0/tag_control_sig_2_0_8[7] ));
    OR2A \data_source_0/tag_data_buf_17_RNO[0]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_17[7]_net_1 ), .Y(
        \data_source_0/tag_data_buf_17_4[0] ));
    NOR2B \data_source_0/tag_control_sig_RNO_18[16]  (.A(
        \data_source_0/N_1245 ), .B(\data_source_0/N_1178 ), .Y(
        \data_source_0/N_1073 ));
    OR3 \data_source_0/tag_control_sig_RNO_13[4]  (.A(
        \data_source_0/N_1163 ), .B(\data_source_0/N_1178 ), .C(
        \data_source_0/N_1160 ), .Y(\data_source_0/N_783 ));
    NOR2B \data_source_0/tag_data_buf_1_RNO[3]  (.A(
        \data_source_0/tag_data_buf_1[2]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_1_4[3] ));
    IOPAD_TRI \output_signal_pad[7]/U0/U0  (.D(
        \output_signal_pad[7]/U0/NET1 ), .E(
        \output_signal_pad[7]/U0/NET2 ), .PAD(output_signal[7]));
    AO1 \data_source_0/tag_control_sig_RNO_5[0]  (.A(
        \data_source_0/N_726 ), .B(\data_source_0/N_1198 ), .C(
        \data_source_0/N_819 ), .Y(
        \data_source_0/tag_control_sig_2_0_8[0] ));
    OR2 \data_source_0/tag_control_sig_RNO_14[8]  (.A(
        \data_source_0/N_1185 ), .B(\data_source_0/N_1175 ), .Y(
        \data_source_0/N_785 ));
    DFN1C0 \data_source_0/counter[11]  (.D(\data_source_0/counter_n11 )
        , .CLK(main_clock_0_clock_out), .CLR(reset_c), .Q(
        \data_source_0/counter[11]_net_1 ));
    NOR3 \main_clock_0/counter_RNIFVEB1[7]  (.A(
        \main_clock_0/counter[6]_net_1 ), .B(
        \main_clock_0/counter[7]_net_1 ), .C(
        \main_clock_0/counter[3]_net_1 ), .Y(
        \main_clock_0/counter14_3 ));
    AND2 AND2_0 (.A(trigger_signal_c), .B(mac_control_signal_c), .Y(
        AND2_0_Y));
    NOR2B \modulator_0/clock_counter_RNIO0O3[2]  (.A(
        \modulator_0/clock_counter_c1 ), .B(
        \modulator_0/clock_counter[2]_net_1 ), .Y(
        \modulator_0/clock_counter_c2 ));
    NOR2B \data_source_0/tag_data_buf_20_RNO[3]  (.A(
        \data_source_0/tag_data_buf_20[2]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_20_4[3] ));
    DFN1E1P0 \data_source_0/tag_data_buf_18[4]  (.D(
        \data_source_0/tag_data_buf_18_4[4] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_18[4]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_11[11]  (.A(
        \data_source_0/N_990 ), .B(\data_source_0/N_997 ), .C(
        \data_source_0/tag_control_sig_2_0_7[11]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_14[11] ));
    OR3 \data_source_0/tag_control_sig_RNO_0[4]  (.A(
        \data_source_0/N_887 ), .B(\data_source_0/N_883 ), .C(
        \data_source_0/tag_control_sig_2_0_3[4] ), .Y(
        \data_source_0/tag_control_sig_2_0_9[4] ));
    DFN1E1P0 \data_source_0/tag_data_buf_12[2]  (.D(
        \data_source_0/tag_data_buf_12_4[2] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_12[2]_net_1 ));
    DFN1P0 \data_source_0/counter[0]  (.D(\data_source_0/counter_n0 ), 
        .CLK(main_clock_0_clock_out), .PRE(reset_c), .Q(
        \data_source_0/counter_i_0[0] ));
    DFN1C0 \data_source_0/data_index_0[7]  (.D(
        \data_source_0/data_index_3[7] ), .CLK(
        modulator_0_output_signal), .CLR(reset_c), .Q(
        \data_source_0/data_index_0[7]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_4[10]  (.A(
        \data_source_0/N_1244 ), .B(\data_source_0/N_1178 ), .Y(
        \data_source_0/N_976 ));
    NOR3C \data_source_0/tag_control_sig_RNO_3[3]  (.A(
        \data_source_0/N_1152 ), .B(\data_source_0/N_704_i ), .C(
        \data_source_0/tag_control_sig_2_0_a20_2_0[3] ), .Y(
        \data_source_0/N_867 ));
    NOR2B \data_source_0/data_index_RNI6H6D[3]  (.A(
        \data_source_0/N_1133 ), .B(
        \data_source_0/data_index[3]_net_1 ), .Y(
        \data_source_0/N_1238 ));
    NOR2B \data_source_0/tag_data_buf_13_RNO[4]  (.A(
        \data_source_0/tag_data_buf_13[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_13_4[4] ));
    NOR2B \data_source_0/tag_control_sig_RNO_14[19]  (.A(
        \data_source_0/N_1205 ), .B(\data_source_0/N_1184 ), .Y(
        \data_source_0/N_1129 ));
    DFN1C0 \modulator_0/counter[1]  (.D(\modulator_0/counter_n1 ), 
        .CLK(main_clock_0_clock_out), .CLR(reset_c), .Q(
        \modulator_0/counter[1]_net_1 ));
    NOR2A \data_source_0/counter_RNIA5EJ[4]  (.A(
        \data_source_0/counter_i_0[4] ), .B(
        \data_source_0/counter[8]_net_1 ), .Y(
        \data_source_0/output_data_1_sqmuxa_i_a3_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_4[0]  (.D(
        \data_source_0/output_data_23[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_4[0]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_21[3]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_3_0[3] ), .B(
        \data_source_0/N_868_1 ), .Y(\data_source_0/N_868 ));
    NOR2B \data_source_0/tag_control_sig_RNO_11[0]  (.A(
        \data_source_0/N_748 ), .B(\data_source_0/N_1183 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_0[0] ));
    DFN1E1C0 \data_source_0/tag_data_buf_6[4]  (.D(
        \data_source_0/tag_data_buf_6_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_6[4]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_5[6]  (.D(
        \data_source_0/tag_data_buf_5_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_5[6]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_2[3]  (.D(
        \data_source_0/tag_data_buf_2_4[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_2[3]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_23[1]  (.A(
        \data_source_0/N_1133 ), .B(\data_source_0/N_1175 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_6_0[1] ));
    AO1 \data_source_0/tag_control_sig_RNO_8[4]  (.A(
        \data_source_0/N_1199 ), .B(\data_source_0/N_1177 ), .C(
        \data_source_0/N_886 ), .Y(
        \data_source_0/tag_control_sig_2_0_4[4] ));
    NOR3C \data_source_0/counter_RNICBKK[6]  (.A(
        \data_source_0/counter_i_0[7] ), .B(
        \data_source_0/counter_i_0[6] ), .C(
        \data_source_0/counter_n9_i_a2_2 ), .Y(
        \data_source_0/counter_n9_i_a2_5 ));
    AX1C \main_clock_0/clock_out_RNO  (.A(\main_clock_0/counter14_3 ), 
        .B(\main_clock_0/counter14_4 ), .C(\main_clock_0/clock_out_i ), 
        .Y(\main_clock_0/clock_out_RNO_net_1 ));
    NOR3B \data_source_0/tag_control_sig_RNO_7[5]  (.A(
        \data_source_0/N_1154 ), .B(\data_source_0/N_1186 ), .C(
        \data_source_0/data_index_0[4]_net_1 ), .Y(
        \data_source_0/N_909 ));
    AO1 \data_source_0/tag_control_sig_RNO_3[14]  (.A(
        \data_source_0/N_1217 ), .B(\data_source_0/N_1162 ), .C(
        \data_source_0/N_886 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[14] ));
    NOR2A \data_source_0/data_index_RNIAL6D[1]  (.A(
        \data_source_0/N_1140 ), .B(
        \data_source_0/data_index[1]_net_1 ), .Y(
        \data_source_0/N_868_1 ));
    OA1 \data_source_0/tag_control_sig_RNO_8[14]  (.A(
        \data_source_0/N_1159 ), .B(\data_source_0/N_1186 ), .C(
        \data_source_0/N_1211 ), .Y(
        \data_source_0/tag_control_sig_2_0_6[14] ));
    OR3 \data_source_0/tag_control_sig_RNO_1[13]  (.A(
        \data_source_0/N_1030 ), .B(\data_source_0/N_1033 ), .C(
        \data_source_0/tag_control_sig_2_0_9[13] ), .Y(
        \data_source_0/tag_control_sig_2_0_14[13] ));
    NOR3C \data_source_0/tag_control_sig_RNO_18[17]  (.A(
        \data_source_0/N_1133 ), .B(\data_source_0/N_1151 ), .C(
        \data_source_0/N_1176 ), .Y(\data_source_0/N_1099 ));
    NOR3C \data_source_0/tag_control_sig_RNO_14[15]  (.A(
        \data_source_0/N_1185 ), .B(\data_source_0/N_1231 ), .C(
        \data_source_0/N_901_1 ), .Y(\data_source_0/N_1057 ));
    DFN1E1C0 \data_source_0/tag_data_buf_19[7]  (.D(
        \data_source_0/tag_data_buf_19_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_19[7]_net_1 ));
    OR2 \data_source_0/tag_control_sig_RNO_17[9]  (.A(
        \data_source_0/N_757 ), .B(\data_source_0/N_1207 ), .Y(
        \data_source_0/N_777 ));
    OR2A \data_source_0/tag_data_buf_8_RNO[3]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_8[2]_net_1 ), .Y(
        \data_source_0/tag_data_buf_8_4[3] ));
    DFN1E1C0 \data_source_0/tag_data_buf_17[2]  (.D(
        \data_source_0/tag_data_buf_17_4[2] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_17[2]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_4[1]  (.A(
        \data_source_0/N_1229 ), .B(\data_source_0/N_1185 ), .Y(
        \data_source_0/N_843 ));
    NOR2B \data_source_0/tag_data_buf_20_RNO[1]  (.A(
        \data_source_0/tag_data_buf_20[0]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_20_4[1] ));
    OR3 \data_source_0/tag_control_sig_RNO_10[1]  (.A(
        \data_source_0/N_832 ), .B(\data_source_0/N_830 ), .C(
        \data_source_0/N_829 ), .Y(
        \data_source_0/tag_control_sig_2_0_9[1] ));
    NOR3C \data_source_0/tag_control_sig_RNO_6[16]  (.A(
        \data_source_0/N_1184 ), .B(\data_source_0/N_668 ), .C(
        \data_source_0/N_1227 ), .Y(\data_source_0/N_1075 ));
    OR3 \data_source_0/tag_control_sig_RNO_10[18]  (.A(
        \data_source_0/N_1109 ), .B(\data_source_0/N_1113 ), .C(
        \data_source_0/tag_control_sig_2_0_6[18] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[18] ));
    NOR2 \modulator_0/counter_RNIPIOV[1]  (.A(
        \modulator_0/counter[0]_net_1 ), .B(
        \modulator_0/counter[1]_net_1 ), .Y(\modulator_0/counter23_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_4[3]  (.D(
        \data_source_0/tag_data_buf_4_4[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_4[3]_net_1 ));
    OR2A \data_source_0/tag_data_buf_15_RNO[2]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_15[1]_net_1 ), .Y(
        \data_source_0/tag_data_buf_15_4[2] ));
    NOR3C \data_source_0/tag_control_sig_RNO_23[9]  (.A(
        \data_source_0/N_1140 ), .B(\data_source_0/N_1154 ), .C(
        \data_source_0/N_1161 ), .Y(\data_source_0/N_970 ));
    NOR3B \data_source_0/tag_control_sig_RNO_21[18]  (.A(
        \data_source_0/N_1191 ), .B(\data_source_0/N_1213 ), .C(
        \data_source_0/data_index[9]_net_1 ), .Y(
        \data_source_0/N_1113 ));
    DFN1E1C0 \data_source_0/output_data[10]  (.D(
        \data_source_0/output_data_23[10] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[10] ));
    NOR2B \data_source_0/tag_data_buf_11_RNO[7]  (.A(
        \data_source_0/tag_data_buf_11[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_11_4[7] ));
    DFN1E1 \data_source_0/tag_control_sig[10]  (.D(
        \data_source_0/tag_control_sig_2[10] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[10] ));
    AO1 \data_source_0/tag_control_sig_RNO_6[11]  (.A(
        \data_source_0/N_1195 ), .B(\data_source_0/N_1162 ), .C(
        \data_source_0/N_1005 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[11] ));
    DFN1C0 \data_source_0/counter[10]  (.D(\data_source_0/counter_n10 )
        , .CLK(main_clock_0_clock_out), .CLR(reset_c), .Q(
        \data_source_0/counter[10]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_20[1]  (.D(
        \data_source_0/tag_data_buf_20_4[1] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_20[1]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_2[13]  (.A(
        \data_source_0/tag_control_sig_2_0_7[13] ), .B(
        \data_source_0/tag_control_sig_2_0_6[13] ), .C(
        \data_source_0/tag_control_sig_2_0_12[13] ), .Y(
        \data_source_0/tag_control_sig_2_0_16[13] ));
    DFN1E1C0 \data_source_0/tag_data_buf_18[6]  (.D(
        \data_source_0/tag_data_buf_18_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_18[6]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_6_RNO[3]  (.A(
        \data_source_0/tag_data_buf_6[2]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_6_4[3] ));
    XAI1 \data_source_0/counter_RNO[2]  (.A(\data_source_0/N_31 ), .B(
        \data_source_0/counter_i_0[2] ), .C(modulator_0_output_signal), 
        .Y(\data_source_0/N_24 ));
    NOR3C \data_source_0/tag_control_sig_RNO_14[13]  (.A(
        \data_source_0/N_1156 ), .B(\data_source_0/N_1155 ), .C(
        \data_source_0/N_1159 ), .Y(\data_source_0/N_1025 ));
    NOR2B \data_source_0/tag_control_sig_RNO_12[1]  (.A(
        \data_source_0/N_1190 ), .B(\data_source_0/N_1179 ), .Y(
        \data_source_0/N_841 ));
    OR2 \data_source_0/data_index_RNI4D731_0[0]  (.A(
        \data_source_0/N_1178 ), .B(\data_source_0/N_1177 ), .Y(
        \data_source_0/N_761 ));
    NOR2B \switching_circuit_0/un90_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[9] ), .B(main_clock_0_clock_out)
        , .Y(\switching_circuit_0/un90_out_signal_switch_0_net_1 ));
    XA1 \modulator_0/clock_counter_RNO[12]  (.A(
        \modulator_0/clock_counter_c11 ), .B(\modulator_0/un6lto12 ), 
        .C(AND2_0_Y), .Y(\modulator_0/clock_counter_n12 ));
    NOR2B \switching_circuit_0/un50_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[5] ), .B(main_clock_0_clock_out)
        , .Y(\switching_circuit_0/un50_out_signal_switch_0_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_4[17]  (.A(
        \data_source_0/N_703_i ), .B(\data_source_0/N_1239 ), .C(
        \data_source_0/tag_control_sig_2_0_a20_2_1[17] ), .Y(
        \data_source_0/N_1089 ));
    OR2 \data_source_0/tag_control_sig_RNO_4[0]  (.A(
        \data_source_0/N_817 ), .B(\data_source_0/N_816 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[0] ));
    NOR3C \data_source_0/tag_control_sig_RNO_19[12]  (.A(
        \data_source_0/N_1136 ), .B(\data_source_0/N_771 ), .C(
        \data_source_0/N_1182 ), .Y(\data_source_0/N_1006 ));
    OR3 \data_source_0/tag_control_sig_RNO_0[10]  (.A(
        \data_source_0/N_980 ), .B(\data_source_0/N_976 ), .C(
        \data_source_0/tag_control_sig_2_0_2[10] ), .Y(
        \data_source_0/tag_control_sig_2_0_8[10] ));
    NOR2B \data_source_0/tag_data_buf_18_RNO[5]  (.A(
        \data_source_0/tag_data_buf_18[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_18_4[5] ));
    CLKIO \reset_pad/U0/U1  (.A(\reset_pad/U0/NET1 ), .Y(reset_c));
    OR3 \data_source_0/tag_control_sig_RNO_10[0]  (.A(
        \data_source_0/N_827 ), .B(
        \data_source_0/tag_control_sig_2_0_6[0] ), .C(
        \data_source_0/tag_control_sig_2_0_5[0] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[0] ));
    DFN1E1 \data_source_0/tag_control_sig[0]  (.D(
        \data_source_0/tag_control_sig_2[0] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[0] ));
    NOR2B \data_source_0/data_index_RNIIF0M_2[6]  (.A(
        \data_source_0/N_1147 ), .B(\data_source_0/N_1152 ), .Y(
        \data_source_0/N_1201 ));
    XA1A \switching_circuit_0/un183_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[18] ), 
        .C(\data_source_0_tag_control_sig[18] ), .Y(
        \switching_circuit_0/un183_out_signal_switch_0_net_1 ));
    MX2 \switching_circuit_0/out_signal_switch_1[14]  (.A(
        \switching_circuit_0/un140_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un143_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[14] ));
    XA1A \data_source_0/tag_control_sig_RNO_22[3]  (.A(
        \data_source_0/data_index[2]_net_1 ), .B(
        \data_source_0/data_index[6]_net_1 ), .C(
        \data_source_0/N_1162 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_3_0[3] ));
    NOR2B \data_source_0/data_index_RNIRO0M_1[7]  (.A(
        \data_source_0/N_1143 ), .B(\data_source_0/N_1132 ), .Y(
        \data_source_0/N_1161 ));
    NOR3B \data_source_0/tag_control_sig_RNO_15[3]  (.A(
        \data_source_0/N_1180 ), .B(\data_source_0/N_1232 ), .C(
        \data_source_0/N_668 ), .Y(\data_source_0/N_869 ));
    DFN1E1 \data_source_0/tag_control_sig[12]  (.D(
        \data_source_0/tag_control_sig_2[12] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[12] ));
    DFN1C0 \data_source_0/data_index[4]  (.D(\data_source_0/I_12 ), 
        .CLK(modulator_0_output_signal), .CLR(reset_c), .Q(
        \data_source_0/data_index[4]_net_1 ));
    NOR2B \data_source_0/data_index_RNIUDQU[1]  (.A(
        \data_source_0/N_1149 ), .B(\data_source_0/N_1161 ), .Y(
        \data_source_0/N_1020_1 ));
    NOR2B \data_source_0/tag_data_buf_13_RNO[1]  (.A(
        \data_source_0/tag_data_buf_13[0]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_13_4[1] ));
    OR2A \data_source_0/tag_data_buf_14_RNO[1]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_14[0]_net_1 ), .Y(
        \data_source_0/tag_data_buf_14_4[1] ));
    OR3 \data_source_0/tag_control_sig_RNO_2[1]  (.A(
        \data_source_0/tag_control_sig_2_0_10[1] ), .B(
        \data_source_0/tag_control_sig_2_0_9[1] ), .C(
        \data_source_0/tag_control_sig_2_0_13[1] ), .Y(
        \data_source_0/tag_control_sig_2_0_16[1] ));
    NOR2B \data_source_0/output_data_RNO[14]  (.A(
        \data_source_0/tag_data_buf_15[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[14] ));
    AO1 \data_source_0/tag_control_sig_RNO_5[2]  (.A(
        \data_source_0/N_1190 ), .B(\data_source_0/N_1173 ), .C(
        \data_source_0/N_856 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[2] ));
    NOR3C \data_source_0/tag_control_sig_RNO_17[7]  (.A(
        \data_source_0/N_1183 ), .B(\data_source_0/N_1144 ), .C(
        \data_source_0/N_748 ), .Y(\data_source_0/N_929 ));
    NOR2 \data_source_0/data_index_RNIH3Q8_0[9]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/data_index[9]_net_1 ), .Y(
        \data_source_0/N_1139 ));
    OR3 \data_source_0/tag_control_sig_RNO[10]  (.A(
        \data_source_0/tag_control_sig_2_0_8[10] ), .B(
        \data_source_0/tag_control_sig_2_0_7[10] ), .C(
        \data_source_0/tag_control_sig_2_0_12[10] ), .Y(
        \data_source_0/tag_control_sig_2[10] ));
    DFN1C0 \data_source_0/counter[15]  (.D(\data_source_0/counter_n15 )
        , .CLK(main_clock_0_clock_out), .CLR(reset_c), .Q(
        \data_source_0/counter[15]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_8_RNO[2]  (.A(
        \data_source_0/tag_data_buf_8[1]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_8_4[2] ));
    NOR2B \data_source_0/tag_control_sig_RNO_6[9]  (.A(
        \data_source_0/N_1216 ), .B(\data_source_0/N_1160 ), .Y(
        \data_source_0/N_962 ));
    XA1A \switching_circuit_0/un23_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[2] ), 
        .C(\data_source_0_tag_control_sig[2] ), .Y(
        \switching_circuit_0/un23_out_signal_switch_0_net_1 ));
    XA1 \modulator_0/clock_counter_RNO[5]  (.A(
        \modulator_0/clock_counter_c4 ), .B(
        \modulator_0/clock_counter[5]_net_1 ), .C(AND2_0_Y), .Y(
        \modulator_0/clock_counter_n5 ));
    OR2 \data_source_0/data_index_0_RNIDE421[7]  (.A(
        \data_source_0/N_1179 ), .B(\data_source_0/N_1160 ), .Y(
        \data_source_0/N_755 ));
    DFN1E1C0 \modulator_0/clock_counter[1]  (.D(
        \modulator_0/clock_counter_n1 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/clock_counter[1]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_5[3]  (.D(
        \data_source_0/tag_data_buf_5_4[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_5[3]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_19_RNO[7]  (.A(
        \data_source_0/tag_data_buf_19[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_19_4[7] ));
    NOR2B \data_source_0/tag_data_buf_8_RNO[5]  (.A(
        \data_source_0/tag_data_buf_8[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_8_4[5] ));
    AOI1D \data_source_0/tag_control_sig_RNO_24[8]  (.A(
        \data_source_0/N_1242 ), .B(\data_source_0/N_1178 ), .C(
        \data_source_0/N_1191 ), .Y(\data_source_0/N_943 ));
    OR3 \data_source_0/tag_control_sig_RNO[12]  (.A(
        \data_source_0/tag_control_sig_2_0_11[12] ), .B(
        \data_source_0/tag_control_sig_2_0_10[12] ), .C(
        \data_source_0/tag_control_sig_2_0_12[12] ), .Y(
        \data_source_0/tag_control_sig_2[12] ));
    NOR3B \data_source_0/tag_control_sig_RNO_3[4]  (.A(
        \data_source_0/N_1154 ), .B(\data_source_0/N_1159 ), .C(
        \data_source_0/data_index[5]_net_1 ), .Y(\data_source_0/N_887 )
        );
    NOR2B \data_source_0/tag_data_buf_6_RNIU95H[7]  (.A(
        \data_source_0/tag_data_buf_6[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[5] ));
    NOR2B \data_source_0/data_index_RNIIF0M_0[6]  (.A(
        \data_source_0/N_1147 ), .B(\data_source_0/N_1149 ), .Y(
        \data_source_0/N_1206 ));
    DFN1C0 \data_source_0/data_index[8]  (.D(\data_source_0/I_23 ), 
        .CLK(modulator_0_output_signal), .CLR(reset_c), .Q(
        \data_source_0/data_index[8]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_9[4]  (.A(
        \data_source_0/N_889 ), .B(\data_source_0/N_895 ), .C(
        \data_source_0/tag_control_sig_2_0_7[4] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[4] ));
    OR3 \data_source_0/tag_control_sig_RNO_8[0]  (.A(
        \data_source_0/N_1223 ), .B(\data_source_0/N_1224 ), .C(
        \data_source_0/N_813 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[0] ));
    AO1 \data_source_0/tag_control_sig_2_0_4[11]  (.A(
        \data_source_0/N_1162 ), .B(\data_source_0/N_1187 ), .C(
        \data_source_0/N_1001 ), .Y(
        \data_source_0/tag_control_sig_2_0_4[11]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_11[12]  (.A(
        \data_source_0/N_1006 ), .B(\data_source_0/N_1013 ), .C(
        \data_source_0/tag_control_sig_2_0_2[12] ), .Y(
        \data_source_0/tag_control_sig_2_0_9[12] ));
    DFN1E1C0 \data_source_0/output_data[3]  (.D(
        \data_source_0/output_data_23[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[3] ));
    NOR2B \modulator_0/clock_counter_RNIPAG7[5]  (.A(
        \modulator_0/clock_counter_c4 ), .B(
        \modulator_0/clock_counter[5]_net_1 ), .Y(
        \modulator_0/clock_counter_c5 ));
    DFN1E1C0 \data_source_0/tag_data_buf_10[5]  (.D(
        \data_source_0/tag_data_buf_10_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_10[5]_net_1 ));
    IOPAD_TRI \output_signal_pad[9]/U0/U0  (.D(
        \output_signal_pad[9]/U0/NET1 ), .E(
        \output_signal_pad[9]/U0/NET2 ), .PAD(output_signal[9]));
    IOPAD_TRI \output_signal_pad[5]/U0/U0  (.D(
        \output_signal_pad[5]/U0/NET1 ), .E(
        \output_signal_pad[5]/U0/NET2 ), .PAD(output_signal[5]));
    OR3 \data_source_0/tag_control_sig_RNO[19]  (.A(
        \data_source_0/tag_control_sig_2_0_11[19] ), .B(
        \data_source_0/tag_control_sig_2_0_10[19] ), .C(
        \data_source_0/tag_control_sig_2_0_12[19] ), .Y(
        \data_source_0/tag_control_sig_2[19] ));
    NOR2B \data_source_0/data_index_RNIIF0M_2[5]  (.A(
        \data_source_0/N_1150 ), .B(\data_source_0/N_1152 ), .Y(
        \data_source_0/N_1204 ));
    AND3 \main_clock_0/un5_counter_1_I_8  (.A(
        \main_clock_0/counter[0]_net_1 ), .B(
        \main_clock_0/counter[1]_net_1 ), .C(
        \main_clock_0/counter[2]_net_1 ), .Y(\main_clock_0/N_6 ));
    DFN1E1C0 \data_source_0/output_data[0]  (.D(
        \data_source_0/output_data_23[0] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[0] ));
    DFN1E1C0 \data_source_0/output_data[4]  (.D(
        \data_source_0/output_data_23[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[4] ));
    XA1 \modulator_0/clock_counter_RNO[2]  (.A(
        \modulator_0/clock_counter[2]_net_1 ), .B(
        \modulator_0/clock_counter_c1 ), .C(AND2_0_Y), .Y(
        \modulator_0/clock_counter_n2 ));
    NOR2B \data_source_0/tag_control_sig_RNO_17[4]  (.A(
        \data_source_0/N_1192 ), .B(\data_source_0/N_1181 ), .Y(
        \data_source_0/N_895 ));
    OR2 \modulator_0/output_signal_RNO_9  (.A(\modulator_0/un6lto12 ), 
        .B(\modulator_0/un6lto11 ), .Y(\modulator_0/un5lto15_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_9[10]  (.A(
        \data_source_0/N_1195 ), .B(\data_source_0/N_1163 ), .C(
        \data_source_0/N_975 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[10] ));
    NOR2B \data_source_0/tag_data_buf_3_RNO[4]  (.A(
        \data_source_0/tag_data_buf_3[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_3_4[4] ));
    OR3 \data_source_0/tag_control_sig_RNO_0[17]  (.A(
        \data_source_0/N_1088 ), .B(\data_source_0/N_1089 ), .C(
        \data_source_0/tag_control_sig_2_0_3[17] ), .Y(
        \data_source_0/tag_control_sig_2_0_10[17] ));
    DFN1E1C0 \data_source_0/tag_data_buf_18[3]  (.D(
        \data_source_0/tag_data_buf_18_4[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_18[3]_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_14[10]  (.A(
        \data_source_0/N_1132 ), .B(\data_source_0/N_1217 ), .C(
        \data_source_0/N_1240 ), .Y(\data_source_0/N_981 ));
    XA1A \data_source_0/data_index_RNI9K6D[1]  (.A(
        \data_source_0/data_index[2]_net_1 ), .B(
        \data_source_0/data_index[6]_net_1 ), .C(
        \data_source_0/data_index[1]_net_1 ), .Y(
        \data_source_0/N_1233 ));
    DFN1E1C0 \data_source_0/tag_data_buf_12[6]  (.D(
        \data_source_0/tag_data_buf_12_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_12[6]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_14[0]  (.D(
        \data_source_0/output_data_23[13] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_14[0]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_3[5]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_1_1[5] ), .B(
        \data_source_0/tag_control_sig_2_0_a20_1_0[5] ), .C(
        \data_source_0/N_900 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[5] ));
    AO1 \data_source_0/tag_control_sig_RNO_21[12]  (.A(
        \data_source_0/N_1213 ), .B(\data_source_0/N_1207 ), .C(
        \data_source_0/N_1010 ), .Y(
        \data_source_0/tag_control_sig_2_0_2[12] ));
    NOR2B \data_source_0/data_index_RNIIMJH[0]  (.A(
        \data_source_0/N_1138 ), .B(\data_source_0/N_1144 ), .Y(
        \data_source_0/N_1162 ));
    NOR3C \data_source_0/tag_control_sig_RNO_4[18]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_2_0[18] ), .B(
        \data_source_0/data_index[3]_net_1 ), .C(
        \data_source_0/tag_control_sig_2_0_a20_2_1[18] ), .Y(
        \data_source_0/N_1105 ));
    NOR3B \data_source_0/tag_control_sig_RNO_21[15]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/data_index[0]_net_1 ), .C(
        \data_source_0/data_index_0[7]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_8_0[15] ));
    NOR2B \data_source_0/data_index_RNIIMJH_0[7]  (.A(
        \data_source_0/N_1145 ), .B(\data_source_0/N_1132 ), .Y(
        \data_source_0/N_1177 ));
    DFN1P0 \data_source_0/counter[7]  (.D(\data_source_0/N_14 ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .Q(
        \data_source_0/counter_i_0[7] ));
    AO1 \data_source_0/tag_control_sig_RNO_5[10]  (.A(
        \data_source_0/N_1196 ), .B(\data_source_0/N_1180 ), .C(
        \data_source_0/N_984 ), .Y(
        \data_source_0/tag_control_sig_2_0_2[10] ));
    NOR2B \data_source_0/counter_RNIE3O01[13]  (.A(
        \data_source_0/counter_n9_i_a2_6 ), .B(
        \data_source_0/counter_n9_i_a2_5 ), .Y(\data_source_0/N_87 ));
    OR2A \data_source_0/tag_data_buf_17_RNO[4]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_17[3]_net_1 ), .Y(
        \data_source_0/tag_data_buf_17_4[4] ));
    NOR2B \data_source_0/data_index_RNIU6731_1[9]  (.A(
        \data_source_0/N_1201 ), .B(\data_source_0/N_1159 ), .Y(
        \data_source_0/N_883 ));
    NOR2B \data_source_0/data_index_RNI46K71_1[2]  (.A(
        \data_source_0/N_1202 ), .B(\data_source_0/N_1174 ), .Y(
        \data_source_0/N_816 ));
    DFN1E1P0 \data_source_0/tag_data_buf_13[0]  (.D(
        \data_source_0/tag_data_buf_13_4[0] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_13[0]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_2[3]  (.A(
        \data_source_0/tag_control_sig_2_0_8[3] ), .B(
        \data_source_0/tag_control_sig_2_0_7[3] ), .C(
        \data_source_0/tag_control_sig_2_0_11[3] ), .Y(
        \data_source_0/tag_control_sig_2_0_14[3] ));
    NOR3C \data_source_0/tag_control_sig_RNO_20[1]  (.A(
        \data_source_0/tag_control_sig_1_3[649] ), .B(
        \data_source_0/N_1148 ), .C(\data_source_0/N_1163 ), .Y(
        \data_source_0/N_848 ));
    MX2 \switching_circuit_0/out_signal_switch_1[19]  (.A(
        \switching_circuit_0/un190_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un193_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[19] ));
    AO1 \data_source_0/tag_control_sig_RNO_7[8]  (.A(
        \data_source_0/N_785 ), .B(\data_source_0/N_1199 ), .C(
        \data_source_0/N_952 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[8] ));
    NOR2B \data_source_0/tag_control_sig_RNO_22[10]  (.A(
        \data_source_0/N_1196 ), .B(\data_source_0/N_1186 ), .Y(
        \data_source_0/N_985 ));
    NOR2B \modulator_0/clock_counter_RNIPVCH1[13]  (.A(
        \modulator_0/clock_counter_c12 ), .B(
        \modulator_0/clock_counter[13]_net_1 ), .Y(
        \modulator_0/clock_counter_c13 ));
    XA1A \switching_circuit_0/un123_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[12] ), 
        .C(\data_source_0_tag_control_sig[12] ), .Y(
        \switching_circuit_0/un123_out_signal_switch_0_net_1 ));
    XAI1 \data_source_0/counter_RNO[7]  (.A(\data_source_0/N_36 ), .B(
        \data_source_0/counter_i_0[7] ), .C(modulator_0_output_signal), 
        .Y(\data_source_0/N_14 ));
    OR3 \data_source_0/tag_control_sig_RNO_10[16]  (.A(
        \data_source_0/N_921 ), .B(\data_source_0/N_1218 ), .C(
        \data_source_0/N_1081 ), .Y(
        \data_source_0/tag_control_sig_2_0_4[16] ));
    DFN1E1C0 \data_source_0/tag_data_buf_13[1]  (.D(
        \data_source_0/tag_data_buf_13_4[1] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_13[1]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_2_RNIQTOS[7]  (.A(
        \data_source_0/tag_data_buf_2[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[1] ));
    XA1A \switching_circuit_0/un103_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[10] ), 
        .C(\data_source_0_tag_control_sig[10] ), .Y(
        \switching_circuit_0/un103_out_signal_switch_0_net_1 ));
    DFN1E1P0 \data_source_0/tag_data_buf_12[3]  (.D(
        \data_source_0/tag_data_buf_12_4[3] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_12[3]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_4[5]  (.A(
        \data_source_0/N_1197 ), .B(\data_source_0/N_1193 ), .Y(
        \data_source_0/N_910 ));
    NOR2B \data_source_0/tag_control_sig_RNO_3[1]  (.A(
        \data_source_0/N_1188 ), .B(\data_source_0/N_1174 ), .Y(
        \data_source_0/N_844 ));
    OA1 \data_source_0/tag_control_sig_RNO_12[19]  (.A(
        \data_source_0/N_1123_1 ), .B(
        \data_source_0/tag_control_sig_2_0_46_tz_0 ), .C(
        \data_source_0/N_1173 ), .Y(
        \data_source_0/tag_control_sig_RNO_12[19]_net_1 ));
    NOR2B \data_source_0/data_index_RNI46K71[1]  (.A(
        \data_source_0/N_1189 ), .B(\data_source_0/N_1174 ), .Y(
        \data_source_0/N_822 ));
    IOTRI_OB_EB \output_signal_pad[7]/U0/U1  (.D(\output_signal_c[7] ), 
        .E(VCC), .DOUT(\output_signal_pad[7]/U0/NET1 ), .EOUT(
        \output_signal_pad[7]/U0/NET2 ));
    AO1 \data_source_0/tag_control_sig_RNO_22[1]  (.A(
        \data_source_0/N_1200 ), .B(\data_source_0/N_1184 ), .C(
        \data_source_0/N_846 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[1] ));
    OA1 \data_source_0/tag_control_sig_RNO_17[0]  (.A(
        \data_source_0/N_1210 ), .B(\data_source_0/N_1225 ), .C(
        \data_source_0/N_1163 ), .Y(
        \data_source_0/tag_control_sig_2_0_6[0] ));
    NOR2B \switching_circuit_0/un70_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[7] ), .B(main_clock_0_clock_out)
        , .Y(\switching_circuit_0/un70_out_signal_switch_0_net_1 ));
    NOR2B \switching_circuit_0/un140_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[14] ), .B(
        main_clock_0_clock_out), .Y(
        \switching_circuit_0/un140_out_signal_switch_0_net_1 ));
    IOTRI_OB_EB \output_signal_pad[12]/U0/U1  (.D(
        \output_signal_c[12] ), .E(VCC), .DOUT(
        \output_signal_pad[12]/U0/NET1 ), .EOUT(
        \output_signal_pad[12]/U0/NET2 ));
    DFN1E1 \data_source_0/tag_control_sig[14]  (.D(
        \data_source_0/tag_control_sig_2[14] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[14] ));
    OR3 \data_source_0/tag_control_sig_RNO_1[15]  (.A(
        \data_source_0/N_1064 ), .B(\data_source_0/N_1071 ), .C(
        \data_source_0/tag_control_sig_2_0_8[15] ), .Y(
        \data_source_0/tag_control_sig_2_0_13[15] ));
    NOR2B \data_source_0/tag_control_sig_RNO_13[19]  (.A(
        \data_source_0/N_1135 ), .B(\data_source_0/N_1144 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_0_0[19] ));
    DFN1E1C0 \data_source_0/tag_data_buf_1[2]  (.D(
        \data_source_0/tag_data_buf_1_4[2] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_1[2]_net_1 ));
    DFN1E1P0 \data_source_0/tag_data_buf_11[0]  (.D(
        \data_source_0/tag_data_buf_11_4[0] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_11[0]_net_1 ));
    NOR2B \data_source_0/data_index_RNI46K71[2]  (.A(
        \data_source_0/N_1217 ), .B(\data_source_0/N_1174 ), .Y(
        \data_source_0/N_873 ));
    OR3 \data_source_0/tag_control_sig_RNO_1[0]  (.A(
        \data_source_0/N_811 ), .B(\data_source_0/N_825 ), .C(
        \data_source_0/tag_control_sig_2_0_7[0] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[0] ));
    OA1 \data_source_0/tag_control_sig_RNO_13[6]  (.A(
        \data_source_0/N_1155 ), .B(\data_source_0/N_1171 ), .C(
        \data_source_0/N_1140 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_1_0[6] ));
    DFN1C0 \data_source_0/data_index[9]  (.D(
        \data_source_0/data_index_3[9] ), .CLK(
        modulator_0_output_signal), .CLR(reset_c), .Q(
        \data_source_0/data_index[9]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_1[3]  (.D(
        \data_source_0/tag_data_buf_1_4[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_1[3]_net_1 ));
    NOR3B \data_source_0/tag_control_sig_RNO_20[0]  (.A(
        \data_source_0/N_1175 ), .B(\data_source_0/N_1136 ), .C(
        \data_source_0/N_759 ), .Y(\data_source_0/N_818 ));
    DFN1E1C0 \data_source_0/tag_data_buf_20[3]  (.D(
        \data_source_0/tag_data_buf_20_4[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_20[3]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_4[3]  (.A(
        \data_source_0/N_1193 ), .B(\data_source_0/N_1190 ), .Y(
        \data_source_0/N_876 ));
    NOR2B \data_source_0/tag_data_buf_3_RNO[6]  (.A(
        \data_source_0/tag_data_buf_3[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_3_4[6] ));
    OR3 \data_source_0/tag_control_sig_RNO_9[17]  (.A(
        \data_source_0/N_1100 ), .B(\data_source_0/N_1099 ), .C(
        \data_source_0/N_1098 ), .Y(
        \data_source_0/tag_control_sig_2_0_8[17] ));
    NOR2B \data_source_0/data_index_RNI46K71_0[2]  (.A(
        \data_source_0/N_1217 ), .B(\data_source_0/N_1181 ), .Y(
        \data_source_0/N_856 ));
    XA1A \switching_circuit_0/un33_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[3] ), 
        .C(\data_source_0_tag_control_sig[3] ), .Y(
        \switching_circuit_0/un33_out_signal_switch_0_net_1 ));
    NOR2B \modulator_0/counter_RNISLOV[4]  (.A(
        \modulator_0/counter[4]_net_1 ), .B(
        \modulator_0/counter[0]_net_1 ), .Y(\modulator_0/counter19_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_12[15]  (.A(
        \data_source_0/N_1226 ), .B(\data_source_0/N_1162 ), .Y(
        \data_source_0/N_1058 ));
    NOR2B \data_source_0/tag_data_buf_15_RNO[4]  (.A(
        \data_source_0/tag_data_buf_15[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_15_4[4] ));
    OR3 \data_source_0/tag_control_sig_RNO_8[6]  (.A(
        \data_source_0/N_817 ), .B(\data_source_0/N_903 ), .C(
        \data_source_0/tag_control_sig_2_0_0[6] ), .Y(
        \data_source_0/tag_control_sig_2_0_9[6] ));
    DFN1C0 \data_source_0/data_index[3]  (.D(
        \data_source_0/data_index_3[3] ), .CLK(
        modulator_0_output_signal), .CLR(reset_c), .Q(
        \data_source_0/data_index[3]_net_1 ));
    DFN1E1C0 \modulator_0/clock_counter[15]  (.D(
        \modulator_0/clock_counter_n15 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/clock_counter[15]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_13_RNO[7]  (.A(
        \data_source_0/tag_data_buf_13[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_13_4[7] ));
    DFN1E1P0 \data_source_0/tag_data_buf_1[0]  (.D(
        \data_source_0/tag_data_buf_1_4[0] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_1[0]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_2[15]  (.A(
        \data_source_0/tag_control_sig_2_0_4[15]_net_1 ), .B(
        \data_source_0/tag_control_sig_2_0_3[15] ), .C(
        \data_source_0/tag_control_sig_2_0_12[15] ), .Y(
        \data_source_0/tag_control_sig_2_0_15[15] ));
    NOR2B \data_source_0/tag_control_sig_RNO_13[15]  (.A(
        \data_source_0/N_1207 ), .B(\data_source_0/N_1174 ), .Y(
        \data_source_0/N_1068 ));
    NOR2B \data_source_0/tag_data_buf_7_RNO[6]  (.A(
        \data_source_0/tag_data_buf_7[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_7_4[6] ));
    NOR2B \data_source_0/tag_data_buf_12_RNIBQSK[7]  (.A(
        \data_source_0/tag_data_buf_12[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[11] ));
    IOTRI_OB_EB \output_signal_pad[15]/U0/U1  (.D(
        \output_signal_c[15] ), .E(VCC), .DOUT(
        \output_signal_pad[15]/U0/NET1 ), .EOUT(
        \output_signal_pad[15]/U0/NET2 ));
    OR3 \data_source_0/tag_control_sig_RNO_0[18]  (.A(
        \data_source_0/N_1111 ), .B(\data_source_0/N_1105 ), .C(
        \data_source_0/tag_control_sig_2_0_3[18] ), .Y(
        \data_source_0/tag_control_sig_2_0_10[18] ));
    XA1A \switching_circuit_0/un163_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[16] ), 
        .C(\data_source_0_tag_control_sig[16] ), .Y(
        \switching_circuit_0/un163_out_signal_switch_0_net_1 ));
    XOR2 \main_clock_0/un5_counter_1_I_17  (.A(\main_clock_0/N_3 ), .B(
        \main_clock_0/counter[6]_net_1 ), .Y(\main_clock_0/I_17_0 ));
    NOR2B \data_source_0/tag_control_sig_RNO_12[9]  (.A(
        \data_source_0/N_1234 ), .B(\data_source_0/N_1144 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_2_0[9] ));
    AO1 \data_source_0/tag_control_sig_RNO_5[17]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_0_0[17] ), .B(
        \data_source_0/N_748 ), .C(\data_source_0/N_1086 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[17] ));
    DFN1E1C0 \data_source_0/tag_data_buf_2[5]  (.D(
        \data_source_0/tag_data_buf_2_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_2[5]_net_1 ));
    IOPAD_IN \clock_pad/U0/U0  (.PAD(clock), .Y(\clock_pad/U0/NET1 ));
    AO1 \data_source_0/tag_control_sig_RNO_10[17]  (.A(
        \data_source_0/N_1213 ), .B(\data_source_0/N_1205 ), .C(
        \data_source_0/N_1097 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[17] ));
    MX2 \switching_circuit_0/out_signal_switch_1[7]  (.A(
        \switching_circuit_0/un70_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un73_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[7] ));
    AND2 \data_source_0/un3_data_index_I_21  (.A(
        \data_source_0/data_index[6]_net_1 ), .B(
        \data_source_0/data_index[7]_net_1 ), .Y(
        \data_source_0/DWACT_FINC_E[3] ));
    OA1 \data_source_0/tag_control_sig_RNO_18[9]  (.A(
        \data_source_0/N_1187 ), .B(\data_source_0/N_1201 ), .C(
        \data_source_0/N_1198 ), .Y(\data_source_0/N_957 ));
    NOR2 \data_source_0/counter_RNI1561[10]  (.A(
        \data_source_0/counter[11]_net_1 ), .B(
        \data_source_0/counter[10]_net_1 ), .Y(
        \data_source_0/counter_n9_i_a2_2 ));
    NOR2A \modulator_0/counter_RNIUNOV[5]  (.A(
        \modulator_0/counter[5]_net_1 ), .B(
        \modulator_0/counter[1]_net_1 ), .Y(\modulator_0/counter19_0 ));
    AOI1D \data_source_0/tag_control_sig_RNO_12[13]  (.A(
        \data_source_0/N_1158 ), .B(\data_source_0/N_1156 ), .C(
        \data_source_0/N_1020_1 ), .Y(\data_source_0/N_1020 ));
    OR3 \data_source_0/tag_control_sig_RNO_0[5]  (.A(
        \data_source_0/tag_control_sig_2_0_0[5] ), .B(
        \data_source_0/N_910 ), .C(
        \data_source_0/tag_control_sig_2_0_7[5] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[5] ));
    NOR2B \modulator_0/output_signal_RNO_11  (.A(\modulator_0/un5lto6 )
        , .B(\modulator_0/clock_counter[5]_net_1 ), .Y(
        \modulator_0/un6lto6_0 ));
    DFN1P0 \data_source_0/data_index[0]  (.D(\data_source_0/I_4 ), 
        .CLK(modulator_0_output_signal), .PRE(reset_c), .Q(
        \data_source_0/data_index[0]_net_1 ));
    NOR2B \modulator_0/clock_counter_RNI2305[3]  (.A(
        \modulator_0/clock_counter_c2 ), .B(
        \modulator_0/clock_counter[3]_net_1 ), .Y(
        \modulator_0/clock_counter_c3 ));
    AOI1D \data_source_0/tag_control_sig_RNO_16[19]  (.A(
        \data_source_0/N_1186 ), .B(\data_source_0/N_1182 ), .C(
        \data_source_0/N_1215 ), .Y(\data_source_0/N_1117 ));
    NOR2B \data_source_0/data_index_RNID81C1[3]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_3_0[9] ), .B(
        \data_source_0/N_853_2 ), .Y(\data_source_0/N_1056 ));
    NOR2B \data_source_0/output_data_RNO[12]  (.A(
        \data_source_0/tag_data_buf_13[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[12] ));
    DFN1E1C0 \data_source_0/tag_data_buf_3[6]  (.D(
        \data_source_0/tag_data_buf_3_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_3[6]_net_1 ));
    DFN1E1P0 \data_source_0/tag_data_buf_15[3]  (.D(
        \data_source_0/tag_data_buf_15_4[3] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_15[3]_net_1 ));
    NOR2A \data_source_0/data_index_RNI1JP8[0]  (.A(
        \data_source_0/data_index[0]_net_1 ), .B(
        \data_source_0/data_index[1]_net_1 ), .Y(
        \data_source_0/tag_control_sig_1_649_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_13[13]  (.A(
        \data_source_0/N_1216 ), .B(\data_source_0/N_1176 ), .Y(
        \data_source_0/N_1035 ));
    AO1 \data_source_0/tag_control_sig_RNO_18[7]  (.A(
        \data_source_0/N_1206 ), .B(\data_source_0/N_1179 ), .C(
        \data_source_0/N_819 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[7] ));
    NOR2B \data_source_0/tag_data_buf_5_RNO[5]  (.A(
        \data_source_0/tag_data_buf_5[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_5_4[5] ));
    DFN1E1C0 \data_source_0/tag_data_buf_15[6]  (.D(
        \data_source_0/tag_data_buf_15_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_15[6]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_11_RNO[4]  (.A(
        \data_source_0/tag_data_buf_11[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_11_4[4] ));
    DFN1E1C0 \modulator_0/clock_counter[5]  (.D(
        \modulator_0/clock_counter_n5 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/clock_counter[5]_net_1 ));
    NOR3A \main_clock_0/counter_RNI0BUP1[2]  (.A(
        \main_clock_0/counter14_2 ), .B(
        \main_clock_0/counter[2]_net_1 ), .C(
        \main_clock_0/counter[5]_net_1 ), .Y(
        \main_clock_0/counter14_4 ));
    NOR2B \data_source_0/tag_data_buf_2_RNO[7]  (.A(
        \data_source_0/tag_data_buf_2[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_2_4[7] ));
    DFN1E1P0 \data_source_0/tag_data_buf_13[2]  (.D(
        \data_source_0/tag_data_buf_13_4[2] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_13[2]_net_1 ));
    AX1C \modulator_0/counter_RNO_0[4]  (.A(
        \modulator_0/counter[3]_net_1 ), .B(\modulator_0/counter_c2 ), 
        .C(\modulator_0/counter[4]_net_1 ), .Y(
        \modulator_0/counter_n4_tz ));
    DFN1E1P0 \data_source_0/tag_data_buf_16[4]  (.D(
        \data_source_0/tag_data_buf_16_4[4] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_16[4]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_16[15]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_8_0[15] ), .B(
        \data_source_0/N_1183 ), .Y(\data_source_0/N_1063 ));
    NOR2B \data_source_0/data_index_RNIIF0M[6]  (.A(
        \data_source_0/N_1147 ), .B(\data_source_0/N_1133 ), .Y(
        \data_source_0/N_1200 ));
    NOR2B \data_source_0/data_index_RNI46K71[5]  (.A(
        \data_source_0/N_1191 ), .B(\data_source_0/N_1184 ), .Y(
        \data_source_0/N_1224 ));
    MX2 \switching_circuit_0/out_signal_switch_1[8]  (.A(
        \switching_circuit_0/un80_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un83_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[8] ));
    OR2A \data_source_0/tag_data_buf_7_RNO[2]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_7[1]_net_1 ), .Y(
        \data_source_0/tag_data_buf_7_4[2] ));
    MX2 \switching_circuit_0/out_signal_switch_1[12]  (.A(
        \switching_circuit_0/un120_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un123_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[12] ));
    IOPAD_TRI \output_signal_pad[11]/U0/U0  (.D(
        \output_signal_pad[11]/U0/NET1 ), .E(
        \output_signal_pad[11]/U0/NET2 ), .PAD(output_signal[11]));
    OR2A \data_source_0/tag_data_buf_15_RNO[0]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_15[7]_net_1 ), .Y(
        \data_source_0/tag_data_buf_15_4[0] ));
    NOR3C \data_source_0/tag_control_sig_RNO_14[4]  (.A(
        \data_source_0/N_1140 ), .B(\data_source_0/N_1149 ), .C(
        \data_source_0/N_1162 ), .Y(\data_source_0/N_888 ));
    OR3 \data_source_0/tag_control_sig_RNO_11[2]  (.A(
        \data_source_0/tag_control_sig_RNO_13[2]_net_1 ), .B(
        \data_source_0/N_851 ), .C(
        \data_source_0/tag_control_sig_2_0_3[2] ), .Y(
        \data_source_0/tag_control_sig_2_0_10[2] ));
    NOR2B \switching_circuit_0/un130_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[13] ), .B(
        main_clock_0_clock_out), .Y(
        \switching_circuit_0/un130_out_signal_switch_0_net_1 ));
    ULSICC_INT INT_ULSICC_INSTANCE_0 (.USTDBY(GND), .LPENA(GND));
    OR2A \data_source_0/counter_RNI3B613[9]  (.A(
        \data_source_0/counter[9]_net_1 ), .B(\data_source_0/N_38 ), 
        .Y(\data_source_0/N_39 ));
    DFN1C0 \modulator_0/counter[3]  (.D(\modulator_0/counter_n3 ), 
        .CLK(main_clock_0_clock_out), .CLR(reset_c), .Q(
        \modulator_0/counter[3]_net_1 ));
    OR2 \data_source_0/data_index_RNIUDQU[9]  (.A(
        \data_source_0/N_1173 ), .B(\data_source_0/N_1159 ), .Y(
        \data_source_0/N_758 ));
    NOR2B \data_source_0/data_index_RNI3LP8[1]  (.A(
        \data_source_0/data_index[1]_net_1 ), .B(
        \data_source_0/data_index[2]_net_1 ), .Y(
        \data_source_0/N_1133 ));
    DFN1E1C0 \data_source_0/tag_data_buf_4[6]  (.D(
        \data_source_0/tag_data_buf_4_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_4[6]_net_1 ));
    OR2A \data_source_0/tag_data_buf_18_RNO[4]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_18[3]_net_1 ), .Y(
        \data_source_0/tag_data_buf_18_4[4] ));
    DFN1P0 \data_source_0/counter[2]  (.D(\data_source_0/N_24 ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .Q(
        \data_source_0/counter_i_0[2] ));
    OA1 \data_source_0/tag_control_sig_RNO_6[6]  (.A(
        \data_source_0/N_1184 ), .B(\data_source_0/N_1198 ), .C(
        \data_source_0/N_1189 ), .Y(\data_source_0/N_914 ));
    AO1 \data_source_0/tag_control_sig_RNO_5[9]  (.A(
        \data_source_0/N_1229 ), .B(\data_source_0/N_1178 ), .C(
        \data_source_0/N_960 ), .Y(
        \data_source_0/tag_control_sig_2_0_8[9] ));
    IOPAD_TRI \output_signal_pad[6]/U0/U0  (.D(
        \output_signal_pad[6]/U0/NET1 ), .E(
        \output_signal_pad[6]/U0/NET2 ), .PAD(output_signal[6]));
    AO1 \data_source_0/tag_control_sig_RNO_9[18]  (.A(
        \data_source_0/N_1211 ), .B(\data_source_0/N_1174 ), .C(
        \data_source_0/N_1102 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[18] ));
    NOR3C \data_source_0/tag_control_sig_RNO_15[11]  (.A(
        \data_source_0/tag_control_sig_1_3[649] ), .B(
        \data_source_0/N_1148 ), .C(\data_source_0/N_1176 ), .Y(
        \data_source_0/N_1005 ));
    OR3 \data_source_0/tag_control_sig_RNO_1[1]  (.A(
        \data_source_0/tag_control_sig_2_0_3[1] ), .B(
        \data_source_0/N_831 ), .C(
        \data_source_0/tag_control_sig_2_0_4[1] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[1] ));
    XOR2 \data_source_0/data_index_RNI7PP8[1]  (.A(
        \data_source_0/data_index[1]_net_1 ), .B(
        \data_source_0/data_index[6]_net_1 ), .Y(
        \data_source_0/N_707_i ));
    NOR2A \data_source_0/data_index_RNIF1Q8_0[7]  (.A(
        \data_source_0/data_index[7]_net_1 ), .B(
        \data_source_0/data_index[8]_net_1 ), .Y(
        \data_source_0/N_1145 ));
    DFN1E1P0 \data_source_0/tag_data_buf_6[1]  (.D(
        \data_source_0/tag_data_buf_6_4[1] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_6[1]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_16[13]  (.A(
        \data_source_0/N_1190 ), .B(\data_source_0/N_1160 ), .Y(
        \data_source_0/N_1024 ));
    NOR2B \data_source_0/tag_data_buf_4_RNO[3]  (.A(
        \data_source_0/tag_data_buf_4[2]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_4_4[3] ));
    NOR2B \data_source_0/tag_control_sig_RNO_7[1]  (.A(
        \data_source_0/N_1183 ), .B(\data_source_0/N_1162 ), .Y(
        \data_source_0/N_831 ));
    DFN1E1C0 \data_source_0/tag_data_buf_6[6]  (.D(
        \data_source_0/tag_data_buf_6_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_6[6]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_16[6]  (.D(
        \data_source_0/tag_data_buf_16_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_16[6]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_11[9]  (.A(
        \data_source_0/N_968 ), .B(\data_source_0/N_967 ), .C(
        \data_source_0/tag_control_sig_2_0_5[9] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[9] ));
    OR3 \data_source_0/tag_control_sig_RNO_10[8]  (.A(
        \data_source_0/N_950 ), .B(\data_source_0/N_951 ), .C(
        \data_source_0/tag_control_sig_2_0_7[8] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[8] ));
    OR3 \data_source_0/tag_control_sig_RNO_2[2]  (.A(
        \data_source_0/tag_control_sig_2_0_2[2] ), .B(
        \data_source_0/tag_control_sig_2_0_1[2] ), .C(
        \data_source_0/tag_control_sig_2_0_10[2] ), .Y(
        \data_source_0/tag_control_sig_2_0_13[2] ));
    AO1 \data_source_0/tag_control_sig_RNO_5[18]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_3_0[18] ), .B(
        \data_source_0/N_1230 ), .C(\data_source_0/N_1114 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[18] ));
    OR2 \data_source_0/counter_RNILOIG1[4]  (.A(
        \data_source_0/counter_i_0[4] ), .B(\data_source_0/N_33 ), .Y(
        \data_source_0/N_34 ));
    OR2A \data_source_0/tag_data_buf_6_RNO[2]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_6[1]_net_1 ), .Y(
        \data_source_0/tag_data_buf_6_4[2] ));
    XOR2 \main_clock_0/un5_counter_1_I_5  (.A(
        \main_clock_0/counter[0]_net_1 ), .B(
        \main_clock_0/counter[1]_net_1 ), .Y(\main_clock_0/I_5_0 ));
    NOR2B \data_source_0/tag_control_sig_RNO_16[6]  (.A(
        \data_source_0/N_1205 ), .B(\data_source_0/N_1185 ), .Y(
        \data_source_0/N_923 ));
    MX2 \switching_circuit_0/out_signal_switch_1[0]  (.A(
        \switching_circuit_0/un1_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un4_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[0] ));
    OR2 \data_source_0/tag_control_sig_RNO_18[3]  (.A(
        \data_source_0/N_1181 ), .B(\data_source_0/N_1159 ), .Y(
        \data_source_0/N_780 ));
    AO1A \data_source_0/tag_control_sig_RNO_13[7]  (.A(
        \data_source_0/data_index_0[4]_net_1 ), .B(
        \data_source_0/N_1148 ), .C(\data_source_0/N_1195 ), .Y(
        \data_source_0/tag_control_sig_2_0_2_tz[7] ));
    IOPAD_TRI \output_signal_pad[2]/U0/U0  (.D(
        \output_signal_pad[2]/U0/NET1 ), .E(
        \output_signal_pad[2]/U0/NET2 ), .PAD(output_signal[2]));
    NOR2A \data_source_0/tag_control_sig_RNO_12[10]  (.A(
        \data_source_0/data_index[5]_net_1 ), .B(
        \data_source_0/data_index[2]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_3_1[10] ));
    DFN1E1C0 \data_source_0/tag_data_buf_10[2]  (.D(
        \data_source_0/tag_data_buf_10_4[2] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_10[2]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_12_RNO[1]  (.A(
        \data_source_0/tag_data_buf_12[0]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_12_4[1] ));
    OR3 \modulator_0/output_signal_RNO_13  (.A(
        \modulator_0/clock_counter[0]_net_1 ), .B(
        \modulator_0/clock_counter[1]_net_1 ), .C(
        \modulator_0/clock_counter[4]_net_1 ), .Y(
        \modulator_0/un6lt4_2 ));
    NOR2B \data_source_0/tag_data_buf_1_RNO[7]  (.A(
        \data_source_0/tag_data_buf_1[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_1_4[7] ));
    XA1 \modulator_0/clock_counter_RNO[11]  (.A(
        \modulator_0/clock_counter_c10 ), .B(\modulator_0/un6lto11 ), 
        .C(AND2_0_Y), .Y(\modulator_0/clock_counter_n11 ));
    DFN1E1P0 \data_source_0/tag_data_buf_6[2]  (.D(
        \data_source_0/tag_data_buf_6_4[2] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_6[2]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_20[0]  (.D(
        \data_source_0/output_data_23[19] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_20[0]_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_14[14]  (.A(
        \data_source_0/N_1140 ), .B(\data_source_0/N_1133 ), .C(
        \data_source_0/N_1173 ), .Y(\data_source_0/N_1046 ));
    NOR2B \data_source_0/tag_data_buf_8_RNO[6]  (.A(
        \data_source_0/tag_data_buf_8[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_8_4[6] ));
    IOTRI_OB_EB \output_signal_pad[9]/U0/U1  (.D(\output_signal_c[9] ), 
        .E(VCC), .DOUT(\output_signal_pad[9]/U0/NET1 ), .EOUT(
        \output_signal_pad[9]/U0/NET2 ));
    IOTRI_OB_EB \output_signal_pad[5]/U0/U1  (.D(\output_signal_c[5] ), 
        .E(VCC), .DOUT(\output_signal_pad[5]/U0/NET1 ), .EOUT(
        \output_signal_pad[5]/U0/NET2 ));
    NOR2B \data_source_0/tag_data_buf_10_RNO[5]  (.A(
        \data_source_0/tag_data_buf_10[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_10_4[5] ));
    OA1 \data_source_0/tag_control_sig_RNO_13[10]  (.A(
        \data_source_0/N_1227 ), .B(\data_source_0/N_1232 ), .C(
        \data_source_0/N_1160 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_3_0[10] ));
    NOR3C \data_source_0/tag_control_sig_RNO_3[10]  (.A(
        \data_source_0/tag_control_sig_1_3[649] ), .B(
        \data_source_0/N_1148 ), .C(\data_source_0/N_1159 ), .Y(
        \data_source_0/N_980 ));
    NOR2B \data_source_0/tag_data_buf_14_RNO[6]  (.A(
        \data_source_0/tag_data_buf_14[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_14_4[6] ));
    AO1 \data_source_0/tag_control_sig_RNO_8[10]  (.A(
        \data_source_0/N_726 ), .B(\data_source_0/N_1181 ), .C(
        \data_source_0/N_982 ), .Y(
        \data_source_0/tag_control_sig_2_0_6[10] ));
    NOR3C \data_source_0/tag_control_sig_RNO_18[5]  (.A(
        \data_source_0/N_1133 ), .B(\data_source_0/N_1151 ), .C(
        \data_source_0/tag_control_sig_2_0_a20_10_0[5] ), .Y(
        \data_source_0/N_908 ));
    OR2 \data_source_0/tag_control_sig_RNO_2[0]  (.A(
        \data_source_0/tag_control_sig_2_0_10[0] ), .B(
        \data_source_0/tag_control_sig_2_0_11[0] ), .Y(
        \data_source_0/tag_control_sig_2_0_14[0] ));
    OR3 \data_source_0/tag_control_sig_RNO_0[9]  (.A(
        \data_source_0/tag_control_sig_2_0_1[9] ), .B(
        \data_source_0/tag_control_sig_2_0_0[9] ), .C(
        \data_source_0/tag_control_sig_2_0_8[9] ), .Y(
        \data_source_0/tag_control_sig_2_0_13[9] ));
    NOR2B \data_source_0/counter_RNIVPDJ_0[1]  (.A(
        \data_source_0/counter_i_0[1] ), .B(
        \data_source_0/counter_i_0[0] ), .Y(\data_source_0/N_90 ));
    NOR2B \data_source_0/tag_data_buf_10_RNO[4]  (.A(
        \data_source_0/tag_data_buf_10[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_10_4[4] ));
    DFN1E1C0 \data_source_0/tag_data_buf_14[5]  (.D(
        \data_source_0/tag_data_buf_14_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_14[5]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_22[9]  (.A(
        \data_source_0/data_index[3]_net_1 ), .B(
        \data_source_0/tag_control_sig_2_0_a20_3_0[9] ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_3_2[9] ));
    XA1A \switching_circuit_0/un43_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[4] ), 
        .C(\data_source_0_tag_control_sig[4] ), .Y(
        \switching_circuit_0/un43_out_signal_switch_0_net_1 ));
    NOR2B \data_source_0/data_index_RNIIMJH[7]  (.A(
        \data_source_0/N_1145 ), .B(\data_source_0/N_1141 ), .Y(
        \data_source_0/N_1181 ));
    NOR2A \data_source_0/data_index_RNIO37D_0[7]  (.A(
        \data_source_0/N_1139 ), .B(
        \data_source_0/data_index[7]_net_1 ), .Y(
        \data_source_0/N_1143 ));
    NOR2B \data_source_0/data_index_RNIIF0M[2]  (.A(
        \data_source_0/N_1157 ), .B(
        \data_source_0/tag_control_sig_1_3[649] ), .Y(
        \data_source_0/N_1210 ));
    NOR2B \data_source_0/data_index_RNIRO0M_3[7]  (.A(
        \data_source_0/N_1139 ), .B(\data_source_0/N_1213 ), .Y(
        \data_source_0/N_1242 ));
    NOR2B \data_source_0/tag_control_sig_RNO_7[13]  (.A(
        \data_source_0/N_1205 ), .B(\data_source_0/N_1179 ), .Y(
        \data_source_0/N_1033 ));
    NOR2B \data_source_0/tag_control_sig_RNO_17[11]  (.A(
        \data_source_0/N_1197 ), .B(\data_source_0/N_1185 ), .Y(
        \data_source_0/N_1000 ));
    AND2 \main_clock_0/un5_counter_1_I_15  (.A(
        \main_clock_0/counter[3]_net_1 ), .B(
        \main_clock_0/counter[4]_net_1 ), .Y(
        \main_clock_0/DWACT_FINC_E[1] ));
    DFN1E1 \data_source_0/tag_control_sig[16]  (.D(
        \data_source_0/tag_control_sig_2[16] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[16] ));
    AND3 \data_source_0/un3_data_index_I_19  (.A(
        \data_source_0/DWACT_FINC_E[0] ), .B(
        \data_source_0/DWACT_FINC_E[2] ), .C(
        \data_source_0/data_index[6]_net_1 ), .Y(\data_source_0/N_4 ));
    NOR2B \data_source_0/tag_control_sig_RNO_19[6]  (.A(
        \data_source_0/N_1202 ), .B(\data_source_0/N_1185 ), .Y(
        \data_source_0/N_924 ));
    DFN1E1C0 \data_source_0/tag_data_buf_3[2]  (.D(
        \data_source_0/tag_data_buf_3_4[2] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_3[2]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_16[2]  (.D(
        \data_source_0/tag_data_buf_16_4[2] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_16[2]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_3[5]  (.D(
        \data_source_0/tag_data_buf_3_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_3[5]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_2[4]  (.A(
        \data_source_0/tag_control_sig_2_0_5[4] ), .B(
        \data_source_0/tag_control_sig_2_0_4[4] ), .C(
        \data_source_0/tag_control_sig_2_0_11[4] ), .Y(
        \data_source_0/tag_control_sig_2_0_13[4] ));
    OR2 \data_source_0/tag_control_sig_RNO_19[19]  (.A(
        \data_source_0/N_1196 ), .B(\data_source_0/N_1183 ), .Y(
        \data_source_0/tag_control_sig_2_0_46_tz_0 ));
    NOR3C \data_source_0/tag_control_sig_RNO_6[7]  (.A(
        \data_source_0/N_1139 ), .B(\data_source_0/N_1132 ), .C(
        \data_source_0/N_1217 ), .Y(\data_source_0/N_936 ));
    OR3A \data_source_0/counter_RNIB5FN2[7]  (.A(
        \data_source_0/counter[8]_net_1 ), .B(\data_source_0/N_36 ), 
        .C(\data_source_0/counter_i_0[7] ), .Y(\data_source_0/N_38 ));
    NOR3C \data_source_0/tag_control_sig_RNO_7[9]  (.A(
        \data_source_0/N_1141 ), .B(\data_source_0/N_1204 ), .C(
        \data_source_0/N_1237 ), .Y(\data_source_0/N_969 ));
    NOR2B \data_source_0/data_index_RNIIF0M[1]  (.A(
        \data_source_0/N_1151 ), .B(\data_source_0/N_1149 ), .Y(
        \data_source_0/N_1229 ));
    IOPAD_TRI \output_signal_pad[1]/U0/U0  (.D(
        \output_signal_pad[1]/U0/NET1 ), .E(
        \output_signal_pad[1]/U0/NET2 ), .PAD(output_signal[1]));
    NOR3C \data_source_0/tag_control_sig_RNO_16[10]  (.A(
        \data_source_0/N_1176 ), .B(\data_source_0/N_707_i ), .C(
        \data_source_0/N_813_1 ), .Y(\data_source_0/N_975 ));
    NOR2B \data_source_0/data_index_RNIU6731_2[9]  (.A(
        \data_source_0/N_1205 ), .B(\data_source_0/N_1159 ), .Y(
        \data_source_0/N_1219 ));
    MX2 \switching_circuit_0/out_signal_switch_1[5]  (.A(
        \switching_circuit_0/un50_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un53_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[5] ));
    OA1B \data_source_0/counter_RNO_2[8]  (.A(\data_source_0/N_36 ), 
        .B(\data_source_0/counter_i_0[7] ), .C(
        \data_source_0/counter[8]_net_1 ), .Y(\data_source_0/N_69 ));
    OR3 \data_source_0/tag_control_sig_RNO_9[1]  (.A(
        \data_source_0/N_833 ), .B(\data_source_0/N_834 ), .C(
        \data_source_0/tag_control_sig_2_0_2[1] ), .Y(
        \data_source_0/tag_control_sig_2_0_10[1] ));
    NOR3B \data_source_0/tag_control_sig_RNO_17[8]  (.A(
        \data_source_0/N_668 ), .B(
        \data_source_0/tag_control_sig_2_0_a20_4_0[8] ), .C(
        \data_source_0/data_index[1]_net_1 ), .Y(\data_source_0/N_947 )
        );
    NOR2B \data_source_0/data_index_RNIBM6D[2]  (.A(
        \data_source_0/tag_control_sig_1_3[649] ), .B(
        \data_source_0/data_index[2]_net_1 ), .Y(
        \data_source_0/N_813_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_1[19]  (.A(
        \data_source_0/N_1056 ), .B(\data_source_0/N_883 ), .C(
        \data_source_0/tag_control_sig_2_0_4[19] ), .Y(
        \data_source_0/tag_control_sig_2_0_10[19] ));
    AO1B \modulator_0/counter_RNIBT613[1]  (.A(
        \modulator_0/counter23_2 ), .B(\modulator_0/counter23_1 ), .C(
        AND2_0_Y), .Y(\modulator_0/clock_countere ));
    DFN1E1C0 \data_source_0/output_data[11]  (.D(
        \data_source_0/output_data_23[11] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[11] ));
    XA1 \modulator_0/clock_counter_RNO[1]  (.A(
        \modulator_0/clock_counter[1]_net_1 ), .B(
        \modulator_0/clock_counter[0]_net_1 ), .C(AND2_0_Y), .Y(
        \modulator_0/clock_counter_n1 ));
    DFN1C0 \main_clock_0/counter[0]  (.D(\main_clock_0/counter_3[0] ), 
        .CLK(GLA), .CLR(reset_c), .Q(\main_clock_0/counter[0]_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_14[5]  (.A(
        \data_source_0/N_701_i ), .B(\data_source_0/N_1177 ), .C(
        \data_source_0/N_1230 ), .Y(\data_source_0/N_900 ));
    OR2A \data_source_0/tag_data_buf_14_RNO[3]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_14[2]_net_1 ), .Y(
        \data_source_0/tag_data_buf_14_4[3] ));
    AO1 \data_source_0/tag_control_sig_RNO_19[15]  (.A(
        \data_source_0/N_1202 ), .B(\data_source_0/N_1186 ), .C(
        \data_source_0/N_1059 ), .Y(
        \data_source_0/tag_control_sig_2_0_6[15] ));
    DFN1E1P0 \data_source_0/tag_data_buf_14[2]  (.D(
        \data_source_0/tag_data_buf_14_4[2] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_14[2]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_3[17]  (.A(
        \data_source_0/N_1245 ), .B(\data_source_0/N_1186 ), .Y(
        \data_source_0/N_1088 ));
    NOR2B \data_source_0/tag_control_sig_RNO_21[10]  (.A(
        \data_source_0/N_1231 ), .B(\data_source_0/N_1193 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_5_0[10] ));
    AND3 \data_source_0/un3_data_index_I_22  (.A(
        \data_source_0/DWACT_FINC_E[0] ), .B(
        \data_source_0/DWACT_FINC_E[2] ), .C(
        \data_source_0/DWACT_FINC_E[3] ), .Y(\data_source_0/N_3 ));
    AO1 \data_source_0/tag_control_sig_RNO_8[17]  (.A(
        \data_source_0/N_1209 ), .B(\data_source_0/N_1175 ), .C(
        \data_source_0/N_1092 ), .Y(
        \data_source_0/tag_control_sig_2_0_2[17] ));
    OR2A \data_source_0/counter_RNO_0[15]  (.A(
        \data_source_0/counter[14]_net_1 ), .B(\data_source_0/N_43 ), 
        .Y(\data_source_0/N_44 ));
    IOPAD_TRI \output_signal_pad[16]/U0/U0  (.D(
        \output_signal_pad[16]/U0/NET1 ), .E(
        \output_signal_pad[16]/U0/NET2 ), .PAD(output_signal[16]));
    DFN1E1C0 \data_source_0/tag_data_buf_13[4]  (.D(
        \data_source_0/tag_data_buf_13_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_13[4]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_8[2]  (.A(
        \data_source_0/N_1199 ), .B(\data_source_0/N_1160 ), .C(
        \data_source_0/N_832 ), .Y(
        \data_source_0/tag_control_sig_2_0_6[2] ));
    NOR2B \data_source_0/data_index_RNICN6D_0[9]  (.A(
        \data_source_0/N_1141 ), .B(
        \data_source_0/data_index[9]_net_1 ), .Y(
        \data_source_0/N_1175 ));
    DFN1C0 \data_source_0/counter[14]  (.D(\data_source_0/counter_n14 )
        , .CLK(main_clock_0_clock_out), .CLR(reset_c), .Q(
        \data_source_0/counter[14]_net_1 ));
    DFN1E1C0 \data_source_0/output_data[12]  (.D(
        \data_source_0/output_data_23[12] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[12] ));
    OR2A \data_source_0/counter_RNI6KV23[12]  (.A(
        \data_source_0/counter[12]_net_1 ), .B(\data_source_0/N_41 ), 
        .Y(\data_source_0/N_42 ));
    AO1 \data_source_0/tag_control_sig_RNO_5[7]  (.A(
        \data_source_0/N_1161 ), .B(
        \data_source_0/tag_control_sig_2_0_2_tz[7] ), .C(
        \data_source_0/N_941 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[7] ));
    NOR2B \modulator_0/clock_counter_RNIUV581[12]  (.A(
        \modulator_0/clock_counter_c11 ), .B(\modulator_0/un6lto12 ), 
        .Y(\modulator_0/clock_counter_c12 ));
    OR3 \data_source_0/tag_control_sig_RNO_1[12]  (.A(
        \data_source_0/N_1018 ), .B(\data_source_0/N_1019 ), .C(
        \data_source_0/tag_control_sig_2_0_4[12] ), .Y(
        \data_source_0/tag_control_sig_2_0_10[12] ));
    AO1 \data_source_0/data_index_RNI4V0C1[2]  (.A(
        \data_source_0/N_1155 ), .B(\data_source_0/N_1156 ), .C(
        \data_source_0/N_1201 ), .Y(\data_source_0/N_726 ));
    XA1 \data_source_0/tag_control_sig_RNO_15[12]  (.A(
        \data_source_0/data_index[2]_net_1 ), .B(
        \data_source_0/data_index[6]_net_1 ), .C(
        \data_source_0/N_1193 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_2_0[12] ));
    OR3 \data_source_0/tag_control_sig_RNO_2[19]  (.A(
        \data_source_0/tag_control_sig_2_0_3[19] ), .B(
        \data_source_0/tag_control_sig_2_0_2[19] ), .C(
        \data_source_0/tag_control_sig_2_0_8[19] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[19] ));
    OR3 \data_source_0/tag_control_sig_RNO[8]  (.A(
        \data_source_0/tag_control_sig_2_0_9[8] ), .B(
        \data_source_0/tag_control_sig_2_0_8[8] ), .C(
        \data_source_0/tag_control_sig_2_0_13[8] ), .Y(
        \data_source_0/tag_control_sig_2[8] ));
    NOR2A \data_source_0/data_index_RNIFQ6D_0[5]  (.A(
        \data_source_0/N_1135 ), .B(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/N_1150 ));
    AO1 \data_source_0/tag_control_sig_RNO_15[2]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_3_0[2] ), .B(
        \data_source_0/N_853_2 ), .C(\data_source_0/N_854 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[2] ));
    DFN1E1 \data_source_0/tag_control_sig[13]  (.D(
        \data_source_0/tag_control_sig_2[13] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[13] ));
    NOR3C \data_source_0/tag_control_sig_RNO_11[19]  (.A(
        \data_source_0/data_index_0[4]_net_1 ), .B(
        \data_source_0/N_1152 ), .C(
        \data_source_0/tag_control_sig_2_0_a20_2_0[19] ), .Y(
        \data_source_0/N_1120 ));
    NOR2B \data_source_0/tag_control_sig_RNO_14[18]  (.A(
        \data_source_0/N_1225 ), .B(\data_source_0/N_1193 ), .Y(
        \data_source_0/N_1114 ));
    DFN1E1C0 \data_source_0/tag_data_buf_11[4]  (.D(
        \data_source_0/tag_data_buf_11_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_11[4]_net_1 ));
    NOR2B \data_source_0/data_index_RNIIF0M_10[6]  (.A(
        \data_source_0/N_1148 ), .B(\data_source_0/N_1156 ), .Y(
        \data_source_0/N_1211 ));
    NOR2B \data_source_0/output_data_RNO[16]  (.A(
        \data_source_0/tag_data_buf_17[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[16] ));
    NOR3B \data_source_0/counter_RNO_1[9]  (.A(\data_source_0/N_87 ), 
        .B(\data_source_0/counter[8]_net_1 ), .C(\data_source_0/N_34 ), 
        .Y(\data_source_0/N_68 ));
    DFN1P0 \data_source_0/counter[4]  (.D(\data_source_0/N_20 ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .Q(
        \data_source_0/counter_i_0[4] ));
    NOR3C \data_source_0/tag_control_sig_RNO_19[13]  (.A(
        \data_source_0/N_1134 ), .B(\data_source_0/N_1152 ), .C(
        \data_source_0/N_1174 ), .Y(\data_source_0/N_1026 ));
    NOR2B \data_source_0/tag_data_buf_15_RNO[6]  (.A(
        \data_source_0/tag_data_buf_15[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_15_4[6] ));
    AO1 \data_source_0/tag_control_sig_RNO_21[9]  (.A(
        \data_source_0/N_1187 ), .B(\data_source_0/N_1186 ), .C(
        \data_source_0/N_970 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[9] ));
    AO1 \data_source_0/tag_control_sig_RNO_20[8]  (.A(
        \data_source_0/N_1204 ), .B(\data_source_0/N_1160 ), .C(
        \data_source_0/N_943 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[8] ));
    AO1A \data_source_0/counter_RNO_0[8]  (.A(\data_source_0/N_34 ), 
        .B(\data_source_0/counter_n8_i_a3_0_0 ), .C(
        \data_source_0/N_69 ), .Y(\data_source_0/counter_n8_i_0 ));
    DFN1E1C0 \data_source_0/tag_data_buf_8[5]  (.D(
        \data_source_0/tag_data_buf_8_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_8[5]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_10[5]  (.A(
        \data_source_0/N_1200 ), .B(\data_source_0/N_1161 ), .C(
        \data_source_0/N_903 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[5] ));
    DFN1E1C0 \modulator_0/clock_counter[10]  (.D(
        \modulator_0/clock_counter_n10 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/un6lto10 ));
    OR2A \data_source_0/tag_data_buf_10_RNO[3]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_10[2]_net_1 ), .Y(
        \data_source_0/tag_data_buf_10_4[3] ));
    OR3 \data_source_0/tag_control_sig_RNO_2[12]  (.A(
        \data_source_0/tag_control_sig_2_0_1[12] ), .B(
        \data_source_0/tag_control_sig_2_0_0[12] ), .C(
        \data_source_0/tag_control_sig_2_0_9[12] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[12] ));
    DFN1E1C0 \data_source_0/tag_data_buf_4[7]  (.D(
        \data_source_0/tag_data_buf_4_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_4[7]_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_11[4]  (.A(
        \data_source_0/tag_control_sig_1_3[649] ), .B(
        \data_source_0/N_1148 ), .C(\data_source_0/N_534_tz ), .Y(
        \data_source_0/tag_control_sig_RNO_11[4]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_10[7]  (.A(
        \data_source_0/N_1207 ), .B(\data_source_0/N_1181 ), .Y(
        \data_source_0/N_939 ));
    NOR3C \data_source_0/tag_control_sig_RNO_23[7]  (.A(
        \data_source_0/N_1133 ), .B(\data_source_0/N_1151 ), .C(
        \data_source_0/N_1193 ), .Y(\data_source_0/N_938 ));
    OR2 \data_source_0/tag_control_sig_RNO_11[15]  (.A(
        \data_source_0/N_1216 ), .B(\data_source_0/N_1195 ), .Y(
        \data_source_0/N_778 ));
    NOR2B \data_source_0/tag_data_buf_4_RNO[5]  (.A(
        \data_source_0/tag_data_buf_4[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_4_4[5] ));
    NOR2B \data_source_0/tag_control_sig_RNO_6[14]  (.A(
        \data_source_0/N_1205 ), .B(\data_source_0/N_1175 ), .Y(
        \data_source_0/N_1044 ));
    NOR3B \data_source_0/counter_RNO[8]  (.A(\data_source_0/N_38 ), .B(
        modulator_0_output_signal), .C(\data_source_0/counter_n8_i_0 ), 
        .Y(\data_source_0/N_12 ));
    AX1C \data_source_0/un3_data_index_I_12  (.A(
        \data_source_0/data_index[3]_net_1 ), .B(
        \data_source_0/DWACT_FINC_E[0] ), .C(
        \data_source_0/data_index_0[4]_net_1 ), .Y(
        \data_source_0/I_12 ));
    NOR3C \data_source_0/tag_control_sig_RNO_3[6]  (.A(
        \data_source_0/N_1159 ), .B(\data_source_0/N_668 ), .C(
        \data_source_0/N_1232 ), .Y(\data_source_0/N_920 ));
    OR3 \data_source_0/tag_control_sig_RNO_1[8]  (.A(
        \data_source_0/N_955 ), .B(\data_source_0/N_953 ), .C(
        \data_source_0/tag_control_sig_2_0_1[8] ), .Y(
        \data_source_0/tag_control_sig_2_0_8[8] ));
    NOR2B \data_source_0/tag_control_sig_RNO_19[0]  (.A(
        \data_source_0/N_1195 ), .B(\data_source_0/N_1173 ), .Y(
        \data_source_0/N_820 ));
    NOR2B \data_source_0/tag_data_buf_18_RNO[3]  (.A(
        \data_source_0/tag_data_buf_18[2]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_18_4[3] ));
    IOTRI_OB_EB \output_signal_pad[14]/U0/U1  (.D(
        \output_signal_c[14] ), .E(VCC), .DOUT(
        \output_signal_pad[14]/U0/NET1 ), .EOUT(
        \output_signal_pad[14]/U0/NET2 ));
    OR2A \data_source_0/tag_data_buf_14_RNO[2]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_14[1]_net_1 ), .Y(
        \data_source_0/tag_data_buf_14_4[2] ));
    DFN1E1C0 \data_source_0/tag_data_buf_2[2]  (.D(
        \data_source_0/tag_data_buf_2_4[2] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_2[2]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_11[13]  (.A(
        \data_source_0/N_1027 ), .B(\data_source_0/N_1026 ), .C(
        \data_source_0/tag_control_sig_2_0_5[13] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[13] ));
    NOR2B \data_source_0/data_index_RNIIF0M_0[5]  (.A(
        \data_source_0/N_1150 ), .B(\data_source_0/N_1136 ), .Y(
        \data_source_0/N_1191 ));
    NOR2B \data_source_0/tag_data_buf_17_RNO[5]  (.A(
        \data_source_0/tag_data_buf_17[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_17_4[5] ));
    OR2 \data_source_0/counter_RNIVPDJ[1]  (.A(
        \data_source_0/counter_i_0[1] ), .B(
        \data_source_0/counter_i_0[0] ), .Y(\data_source_0/N_31 ));
    DFN1E1C0 \modulator_0/clock_counter[4]  (.D(
        \modulator_0/clock_counter_n4 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/clock_counter[4]_net_1 ));
    NOR2A \data_source_0/tag_control_sig_RNO_17[12]  (.A(
        \data_source_0/N_1134 ), .B(
        \data_source_0/data_index[2]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_1_1[12] ));
    DFN1E1C0 \data_source_0/tag_data_buf_12[0]  (.D(
        \data_source_0/output_data_23[11] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_12[0]_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_19[8]  (.A(
        \data_source_0/N_1136 ), .B(\data_source_0/N_1135 ), .C(
        \data_source_0/N_1185 ), .Y(\data_source_0/N_951 ));
    NOR2A \modulator_0/clock_counter_RNO[0]  (.A(AND2_0_Y), .B(
        \modulator_0/clock_counter[0]_net_1 ), .Y(\modulator_0/N_121 ));
    NOR2B \data_source_0/tag_data_buf_5_RNO[7]  (.A(
        \data_source_0/tag_data_buf_5[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_5_4[7] ));
    DFN1E1C0 \data_source_0/tag_data_buf_10[4]  (.D(
        \data_source_0/tag_data_buf_10_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_10[4]_net_1 ));
    AOI1 \main_clock_0/counter_RNO[0]  (.A(\main_clock_0/counter14_4 ), 
        .B(\main_clock_0/counter14_3 ), .C(
        \main_clock_0/counter[0]_net_1 ), .Y(
        \main_clock_0/counter_3[0] ));
    OR3 \data_source_0/tag_control_sig_RNO_1[16]  (.A(
        \data_source_0/N_1075 ), .B(\data_source_0/N_1076 ), .C(
        \data_source_0/tag_control_sig_2_0_1[16] ), .Y(
        \data_source_0/tag_control_sig_2_0_8[16] ));
    OR2A \data_source_0/tag_data_buf_10_RNO[1]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_10[0]_net_1 ), .Y(
        \data_source_0/tag_data_buf_10_4[1] ));
    NOR3B \data_source_0/tag_control_sig_RNO_3[18]  (.A(
        \data_source_0/N_1154 ), .B(\data_source_0/N_1174 ), .C(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/N_1111 ));
    OR3 \data_source_0/tag_control_sig_RNO[14]  (.A(
        \data_source_0/tag_control_sig_2_0_13[14] ), .B(
        \data_source_0/tag_control_sig_2_0_12[14] ), .C(
        \data_source_0/tag_control_sig_2_0_14[14] ), .Y(
        \data_source_0/tag_control_sig_2[14] ));
    NOR2B \data_source_0/output_data_RNO[4]  (.A(
        \data_source_0/tag_data_buf_5[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[4] ));
    NOR3B \data_source_0/tag_control_sig_RNO_16[2]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/N_1134 ), .C(
        \data_source_0/data_index_0[7]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_3_0[2] ));
    NOR2B \data_source_0/data_index_RNIIMJH_2[7]  (.A(
        \data_source_0/N_1144 ), .B(\data_source_0/N_1142 ), .Y(
        \data_source_0/N_1193 ));
    AO1 \data_source_0/tag_control_sig_RNO_8[18]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_1_0[18] ), .B(
        \data_source_0/N_1243 ), .C(
        \data_source_0/tag_control_sig_2_0_0[18] ), .Y(
        \data_source_0/tag_control_sig_2_0_8[18] ));
    XNOR2 \data_source_0/data_index_RNI7PP8[5]  (.A(
        \data_source_0/data_index[5]_net_1 ), .B(
        \data_source_0/data_index[2]_net_1 ), .Y(\data_source_0/N_668 )
        );
    NOR2A \data_source_0/data_index_RNI9K6D_1[6]  (.A(
        \data_source_0/N_1133 ), .B(
        \data_source_0/data_index[6]_net_1 ), .Y(
        \data_source_0/N_1171 ));
    IOPAD_TRI \output_signal_pad[19]/U0/U0  (.D(
        \output_signal_pad[19]/U0/NET1 ), .E(
        \output_signal_pad[19]/U0/NET2 ), .PAD(output_signal[19]));
    OR3 \data_source_0/tag_control_sig_RNO_1[11]  (.A(
        \data_source_0/tag_control_sig_2_0_0[11] ), .B(
        \data_source_0/N_991 ), .C(
        \data_source_0/tag_control_sig_2_0_9[11] ), .Y(
        \data_source_0/tag_control_sig_2_0_15[11] ));
    XAI1 \data_source_0/counter_RNO[1]  (.A(
        \data_source_0/counter_i_0[0] ), .B(
        \data_source_0/counter_i_0[1] ), .C(modulator_0_output_signal), 
        .Y(\data_source_0/N_26 ));
    IOTRI_OB_EB \output_signal_pad[6]/U0/U1  (.D(\output_signal_c[6] ), 
        .E(VCC), .DOUT(\output_signal_pad[6]/U0/NET1 ), .EOUT(
        \output_signal_pad[6]/U0/NET2 ));
    NOR2B \data_source_0/tag_control_sig_RNO_14[7]  (.A(
        \data_source_0/N_1188 ), .B(\data_source_0/N_1163 ), .Y(
        \data_source_0/N_941 ));
    XA1 \modulator_0/counter_RNO[1]  (.A(
        \modulator_0/counter[0]_net_1 ), .B(
        \modulator_0/counter[1]_net_1 ), .C(
        \modulator_0/counter_0_sqmuxa ), .Y(\modulator_0/counter_n1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_17[6]  (.D(
        \data_source_0/tag_data_buf_17_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_17[6]_net_1 ));
    MX2 \switching_circuit_0/out_signal_switch_1[18]  (.A(
        \switching_circuit_0/un180_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un183_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[18] ));
    OR2B \data_source_0/counter_RNO[0]  (.A(
        \data_source_0/counter_i_0[0] ), .B(modulator_0_output_signal), 
        .Y(\data_source_0/counter_n0 ));
    AND2 \data_source_0/tag_control_sig_2_0_a20_6[11]  (.A(
        \data_source_0/N_1160 ), .B(\data_source_0/N_1191 ), .Y(
        \data_source_0/N_994 ));
    NOR2 \modulator_0/counter_RNITMOV[2]  (.A(
        \modulator_0/counter[2]_net_1 ), .B(
        \modulator_0/counter[3]_net_1 ), .Y(\modulator_0/counter19_3 ));
    OR3 \data_source_0/tag_control_sig_RNO_2[16]  (.A(
        \data_source_0/tag_control_sig_2_0_5[16] ), .B(
        \data_source_0/tag_control_sig_2_0_4[16] ), .C(
        \data_source_0/tag_control_sig_2_0_11[16] ), .Y(
        \data_source_0/tag_control_sig_2_0_13[16] ));
    OR3 \data_source_0/tag_control_sig_RNO_19[10]  (.A(
        \data_source_0/N_1220 ), .B(\data_source_0/N_1219 ), .C(
        \data_source_0/N_985 ), .Y(
        \data_source_0/tag_control_sig_2_0_4[10] ));
    XAI1 \data_source_0/counter_RNO[3]  (.A(\data_source_0/N_32 ), .B(
        \data_source_0/counter_i_0[3] ), .C(modulator_0_output_signal), 
        .Y(\data_source_0/N_22 ));
    XA1 \modulator_0/clock_counter_RNO[10]  (.A(
        \modulator_0/clock_counter_c9 ), .B(\modulator_0/un6lto10 ), 
        .C(AND2_0_Y), .Y(\modulator_0/clock_counter_n10 ));
    NOR2B \data_source_0/tag_control_sig_RNO_13[14]  (.A(
        \data_source_0/N_761 ), .B(\data_source_0/N_1199 ), .Y(
        \data_source_0/N_1038 ));
    MX2 \switching_circuit_0/out_signal_switch_1[9]  (.A(
        \switching_circuit_0/un90_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un93_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[9] ));
    OR3 \data_source_0/tag_control_sig_RNO_2[11]  (.A(
        \data_source_0/tag_control_sig_2_0_6[11] ), .B(
        \data_source_0/tag_control_sig_2_0_5[11] ), .C(
        \data_source_0/tag_control_sig_2_0_14[11] ), .Y(
        \data_source_0/tag_control_sig_2_0_17[11] ));
    NOR2B \data_source_0/data_index_0_RNIJ6UA1_0[7]  (.A(
        \data_source_0/N_1198 ), .B(\data_source_0/N_1189 ), .Y(
        \data_source_0/N_1010 ));
    NOR2B \data_source_0/tag_control_sig_RNO_24[5]  (.A(
        \data_source_0/N_1211 ), .B(\data_source_0/N_1178 ), .Y(
        \data_source_0/N_902 ));
    NOR2B \data_source_0/tag_control_sig_RNO_7[15]  (.A(
        \data_source_0/N_1215 ), .B(\data_source_0/N_1163 ), .Y(
        \data_source_0/N_1071 ));
    NOR3C \data_source_0/tag_control_sig_RNO_15[1]  (.A(
        \data_source_0/N_1136 ), .B(\data_source_0/N_1140 ), .C(
        \data_source_0/N_1160 ), .Y(\data_source_0/N_837 ));
    MX2 \switching_circuit_0/out_signal_switch_1[13]  (.A(
        \switching_circuit_0/un130_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un133_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[13] ));
    DFN1E1P0 \data_source_0/tag_data_buf_7[1]  (.D(
        \data_source_0/tag_data_buf_7_4[1] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_7[1]_net_1 ));
    DFN1E1C0 \data_source_0/output_data[14]  (.D(
        \data_source_0/output_data_23[14] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[14] ));
    DFN1C0 \data_source_0/data_index[1]  (.D(
        \data_source_0/data_index_3[1] ), .CLK(
        modulator_0_output_signal), .CLR(reset_c), .Q(
        \data_source_0/data_index[1]_net_1 ));
    OR3 \modulator_0/output_signal_RNO_12  (.A(
        \modulator_0/clock_counter[2]_net_1 ), .B(
        \modulator_0/clock_counter[3]_net_1 ), .C(
        \modulator_0/un6lt4_2 ), .Y(\modulator_0/un6lto4 ));
    DFN1E1C0 \modulator_0/clock_counter[8]  (.D(
        \modulator_0/clock_counter_n8 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/clock_counter[8]_net_1 ));
    IOTRI_OB_EB \output_signal_pad[2]/U0/U1  (.D(\output_signal_c[2] ), 
        .E(VCC), .DOUT(\output_signal_pad[2]/U0/NET1 ), .EOUT(
        \output_signal_pad[2]/U0/NET2 ));
    DFN1E1P0 \data_source_0/tag_data_buf_19[4]  (.D(
        \data_source_0/tag_data_buf_19_4[4] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_19[4]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_3[9]  (.A(
        \data_source_0/N_1245 ), .B(\data_source_0/N_1177 ), .C(
        \data_source_0/N_816 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[9] ));
    DFN1E1P0 \data_source_0/tag_data_buf_7[0]  (.D(
        \data_source_0/tag_data_buf_7_4[0] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_7[0]_net_1 ));
    NOR2B \data_source_0/data_index_RNIIF0M_3[2]  (.A(
        \data_source_0/N_1155 ), .B(
        \data_source_0/tag_control_sig_1_3[649] ), .Y(
        \data_source_0/N_1215 ));
    DFN1E1P0 \data_source_0/tag_data_buf_3[0]  (.D(
        \data_source_0/tag_data_buf_3_4[0] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_3[0]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_11[5]  (.D(
        \data_source_0/tag_data_buf_11_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_11[5]_net_1 ));
    OR2A \data_source_0/tag_data_buf_11_RNO[1]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_11[0]_net_1 ), .Y(
        \data_source_0/tag_data_buf_11_4[1] ));
    NOR3B \data_source_0/data_index_0_RNI1NTK_1[7]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/N_1132 ), .C(
        \data_source_0/data_index_0[7]_net_1 ), .Y(
        \data_source_0/N_1179 ));
    DFN1E1C0 \data_source_0/tag_data_buf_7[3]  (.D(
        \data_source_0/tag_data_buf_7_4[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_7[3]_net_1 ));
    OR2A \data_source_0/tag_data_buf_15_RNO[3]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_15[2]_net_1 ), .Y(
        \data_source_0/tag_data_buf_15_4[3] ));
    OR3 \data_source_0/tag_control_sig_RNO_11[1]  (.A(
        \data_source_0/N_848 ), .B(\data_source_0/N_847 ), .C(
        \data_source_0/tag_control_sig_2_0_7[1] ), .Y(
        \data_source_0/tag_control_sig_2_0_13[1] ));
    AO1 \data_source_0/tag_control_sig_RNO_4[13]  (.A(
        \data_source_0/N_1209 ), .B(\data_source_0/N_1175 ), .C(
        \data_source_0/N_1020 ), .Y(
        \data_source_0/tag_control_sig_2_0_2[13] ));
    NOR2B \data_source_0/tag_control_sig_RNO_16[3]  (.A(
        \data_source_0/N_1020_1 ), .B(\data_source_0/N_1208 ), .Y(
        \data_source_0/N_875 ));
    DFN1P0 \data_source_0/counter[3]  (.D(\data_source_0/N_22 ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .Q(
        \data_source_0/counter_i_0[3] ));
    XOR2 \data_source_0/un3_data_index_I_5  (.A(
        \data_source_0/data_index[0]_net_1 ), .B(
        \data_source_0/data_index[1]_net_1 ), .Y(\data_source_0/I_5 ));
    AX1C \data_source_0/un3_data_index_I_7  (.A(
        \data_source_0/data_index[1]_net_1 ), .B(
        \data_source_0/data_index[0]_net_1 ), .C(
        \data_source_0/data_index[2]_net_1 ), .Y(\data_source_0/I_7 ));
    NOR3B \data_source_0/tag_control_sig_RNO_14[16]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/N_1135 ), .C(
        \data_source_0/data_index_0[7]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_1_0[16] ));
    DFN1E1C0 \data_source_0/tag_data_buf_20[6]  (.D(
        \data_source_0/tag_data_buf_20_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_20[6]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_17[3]  (.A(
        \data_source_0/N_1201 ), .B(\data_source_0/N_1173 ), .C(
        \data_source_0/N_868 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[3] ));
    DFN1E1P0 \data_source_0/tag_data_buf_15[0]  (.D(
        \data_source_0/tag_data_buf_15_4[0] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_15[0]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_11[10]  (.A(
        \data_source_0/N_1190 ), .B(\data_source_0/N_1177 ), .Y(
        \data_source_0/N_984 ));
    AO1 \data_source_0/tag_control_sig_RNO_9[6]  (.A(
        \data_source_0/N_1197 ), .B(\data_source_0/N_1182 ), .C(
        \data_source_0/N_923 ), .Y(
        \data_source_0/tag_control_sig_2_0_8[6] ));
    NOR2B \data_source_0/data_index_RNICGJH[1]  (.A(
        \data_source_0/tag_control_sig_1_3[649] ), .B(
        \data_source_0/N_1136 ), .Y(\data_source_0/N_1239 ));
    OR2 \data_source_0/data_index_RNI7G731[9]  (.A(
        \data_source_0/N_1175 ), .B(\data_source_0/N_1161 ), .Y(
        \data_source_0/N_729 ));
    NOR3C \modulator_0/clock_counter_RNO_0[15]  (.A(AND2_0_Y), .B(
        \modulator_0/clock_counter[14]_net_1 ), .C(
        \modulator_0/clock_counter_c13 ), .Y(\modulator_0/N_89 ));
    NOR3C \data_source_0/data_index_RNIU6731[5]  (.A(
        \data_source_0/N_1133 ), .B(\data_source_0/N_1151 ), .C(
        \data_source_0/N_1160 ), .Y(\data_source_0/N_1223 ));
    NOR2B \data_source_0/tag_control_sig_RNO_21[4]  (.A(
        \data_source_0/N_1206 ), .B(\data_source_0/N_1174 ), .Y(
        \data_source_0/N_894 ));
    OA1A \data_source_0/tag_control_sig_RNO_20[7]  (.A(
        \data_source_0/data_index[3]_net_1 ), .B(
        \data_source_0/data_index[7]_net_1 ), .C(
        \data_source_0/N_1196 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_0[7] ));
    NOR2B \data_source_0/tag_control_sig_RNO_16[14]  (.A(
        \data_source_0/N_1191 ), .B(\data_source_0/N_1163 ), .Y(
        \data_source_0/N_1052 ));
    NOR3B \data_source_0/tag_control_sig_RNO_20[16]  (.A(
        \data_source_0/N_1157 ), .B(
        \data_source_0/data_index[8]_net_1 ), .C(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_2[16] ));
    NOR2B \data_source_0/tag_data_buf_16_RNO[6]  (.A(
        \data_source_0/tag_data_buf_16[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_16_4[6] ));
    DFN1E1P0 \data_source_0/tag_data_buf_11[1]  (.D(
        \data_source_0/tag_data_buf_11_4[1] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_11[1]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_16[3]  (.D(
        \data_source_0/tag_data_buf_16_4[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_16[3]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_3[8]  (.A(
        \data_source_0/N_766 ), .B(\data_source_0/N_1176 ), .Y(
        \data_source_0/N_945 ));
    OR3 \data_source_0/tag_control_sig_RNO_11[5]  (.A(
        \data_source_0/N_897 ), .B(\data_source_0/N_908 ), .C(
        \data_source_0/tag_control_sig_2_0_1[5] ), .Y(
        \data_source_0/tag_control_sig_2_0_9[5] ));
    XOR2 \data_source_0/data_index_RNI5NP8[0]  (.A(
        \data_source_0/data_index[0]_net_1 ), .B(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/N_704_i ));
    NOR2B \data_source_0/data_index_RNI7PP8_0[1]  (.A(
        \data_source_0/data_index[1]_net_1 ), .B(
        \data_source_0/data_index[6]_net_1 ), .Y(
        \data_source_0/N_1231 ));
    IOTRI_OB_EB \output_signal_pad[1]/U0/U1  (.D(\output_signal_c[1] ), 
        .E(VCC), .DOUT(\output_signal_pad[1]/U0/NET1 ), .EOUT(
        \output_signal_pad[1]/U0/NET2 ));
    OR2 \data_source_0/counter_RNIUS042[6]  (.A(\data_source_0/N_35 ), 
        .B(\data_source_0/counter_i_0[6] ), .Y(\data_source_0/N_36 ));
    NOR2B \data_source_0/tag_data_buf_14_RNID03N[7]  (.A(
        \data_source_0/tag_data_buf_14[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[13] ));
    NOR2A \data_source_0/data_index_RNIBM6D_0[4]  (.A(
        \data_source_0/N_1137 ), .B(
        \data_source_0/data_index[4]_net_1 ), .Y(
        \data_source_0/N_1227 ));
    NOR2B \data_source_0/output_data_RNO[0]  (.A(
        \data_source_0/tag_data_buf_1[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[0] ));
    DFN1E1C0 \data_source_0/output_data[6]  (.D(
        \data_source_0/output_data_23[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[6] ));
    XOR2 \data_source_0/un3_data_index_I_17  (.A(\data_source_0/N_5 ), 
        .B(\data_source_0/data_index[6]_net_1 ), .Y(
        \data_source_0/I_17 ));
    NOR2B \modulator_0/clock_counter_RNIB3OL[10]  (.A(
        \modulator_0/clock_counter_c9 ), .B(\modulator_0/un6lto10 ), 
        .Y(\modulator_0/clock_counter_c10 ));
    AO1 \data_source_0/tag_control_sig_RNO_4[8]  (.A(
        \data_source_0/N_800 ), .B(\data_source_0/N_1195 ), .C(
        \data_source_0/N_954 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[8] ));
    NOR2B \data_source_0/tag_control_sig_RNO_12[18]  (.A(
        \data_source_0/N_1144 ), .B(\data_source_0/N_704_i ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_2_1[18] ));
    OR2A \data_source_0/tag_data_buf_7_RNO[1]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_7[0]_net_1 ), .Y(
        \data_source_0/tag_data_buf_7_4[1] ));
    XA1A \switching_circuit_0/un173_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[17] ), 
        .C(\data_source_0_tag_control_sig[17] ), .Y(
        \switching_circuit_0/un173_out_signal_switch_0_net_1 ));
    XA1A \switching_circuit_0/un4_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[0] ), 
        .C(\data_source_0_tag_control_sig[0] ), .Y(
        \switching_circuit_0/un4_out_signal_switch_0_net_1 ));
    NOR2B \data_source_0/tag_data_buf_16_RNO[3]  (.A(
        \data_source_0/tag_data_buf_16[2]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_16_4[3] ));
    NOR2B \data_source_0/tag_data_buf_12_RNO[4]  (.A(
        \data_source_0/tag_data_buf_12[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_12_4[4] ));
    DFN1E1C0 \data_source_0/tag_data_buf_13[7]  (.D(
        \data_source_0/tag_data_buf_13_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_13[7]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_0[1]  (.A(
        \data_source_0/N_844 ), .B(\data_source_0/N_843 ), .C(
        \data_source_0/tag_control_sig_2_0_5[1] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[1] ));
    NOR2B \data_source_0/tag_control_sig_RNO_14[17]  (.A(
        \data_source_0/N_758 ), .B(\data_source_0/N_1189 ), .Y(
        \data_source_0/N_1086 ));
    NOR2B \data_source_0/tag_control_sig_RNO_13[18]  (.A(
        \data_source_0/N_701_i ), .B(\data_source_0/N_1180 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_3_0[18] ));
    AOI1B \data_source_0/data_index_RNO[3]  (.A(
        \data_source_0/tag_control_sig_1_649_6 ), .B(
        \data_source_0/tag_control_sig_1_3[649] ), .C(
        \data_source_0/I_9 ), .Y(\data_source_0/data_index_3[3] ));
    NOR2B \data_source_0/data_index_RNIRO0M_0[7]  (.A(
        \data_source_0/N_1143 ), .B(\data_source_0/N_1142 ), .Y(
        \data_source_0/N_1186 ));
    DFN1E1C0 \modulator_0/clock_counter[7]  (.D(
        \modulator_0/clock_counter_n7 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/clock_counter[7]_net_1 ));
    DFN1E1P0 \data_source_0/tag_data_buf_15[1]  (.D(
        \data_source_0/tag_data_buf_15_4[1] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_15[1]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_6[3]  (.D(
        \data_source_0/tag_data_buf_6_4[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_6[3]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_15[0]  (.A(
        \data_source_0/N_1244 ), .B(\data_source_0/N_1182 ), .C(
        \data_source_0/N_820 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[0] ));
    DFN1E1C0 \data_source_0/tag_data_buf_1[6]  (.D(
        \data_source_0/tag_data_buf_1_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_1[6]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_9[0]  (.A(
        \data_source_0/N_815 ), .B(\data_source_0/N_823 ), .C(
        \data_source_0/tag_control_sig_2_0_3[0] ), .Y(
        \data_source_0/tag_control_sig_2_0_10[0] ));
    OR3 \data_source_0/tag_control_sig_RNO_0[13]  (.A(
        \data_source_0/tag_control_sig_2_0_3[13] ), .B(
        \data_source_0/tag_control_sig_2_0_2[13] ), .C(
        \data_source_0/tag_control_sig_2_0_10[13] ), .Y(
        \data_source_0/tag_control_sig_2_0_15[13] ));
    DFN1E1C0 \data_source_0/tag_data_buf_1[7]  (.D(
        \data_source_0/tag_data_buf_1_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_1[7]_net_1 ));
    NOR2B \data_source_0/data_index_RNIIF0M_0[1]  (.A(
        \data_source_0/N_1151 ), .B(\data_source_0/N_1152 ), .Y(
        \data_source_0/N_1189 ));
    NOR2B \data_source_0/tag_control_sig_RNO_24[7]  (.A(
        \data_source_0/N_707_i ), .B(\data_source_0/N_1177 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_2_0[7] ));
    NOR2B \data_source_0/data_index_RNIU6731_0[9]  (.A(
        \data_source_0/N_1215 ), .B(\data_source_0/N_1175 ), .Y(
        \data_source_0/N_833 ));
    DFN1E1 \data_source_0/tag_control_sig[7]  (.D(
        \data_source_0/tag_control_sig_2[7] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[7] ));
    AO1B \data_source_0/counter_RNIK0AI3[1]  (.A(
        \data_source_0/output_data_1_sqmuxa_i_a3_4 ), .B(
        \data_source_0/N_87 ), .C(modulator_0_output_signal), .Y(
        \data_source_0/counter_RNIK0AI3[1]_net_1 ));
    DFN1P0 \data_source_0/counter[1]  (.D(\data_source_0/N_26 ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .Q(
        \data_source_0/counter_i_0[1] ));
    DFN1E1C0 \data_source_0/tag_data_buf_12[4]  (.D(
        \data_source_0/tag_data_buf_12_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_12[4]_net_1 ));
    NOR2B \modulator_0/counter_RNO[2]  (.A(
        \modulator_0/counter_0_sqmuxa ), .B(
        \modulator_0/counter_n2_tz ), .Y(\modulator_0/counter_n2 ));
    AO1A \data_source_0/counter_RNO_0[9]  (.A(
        \data_source_0/counter[9]_net_1 ), .B(\data_source_0/N_38 ), 
        .C(\data_source_0/N_68 ), .Y(\data_source_0/counter_n9_i_0 ));
    NOR3B \data_source_0/counter_RNO[9]  (.A(\data_source_0/N_39 ), .B(
        modulator_0_output_signal), .C(\data_source_0/counter_n9_i_0 ), 
        .Y(\data_source_0/N_10 ));
    NOR3C \data_source_0/tag_control_sig_RNO_11[7]  (.A(
        \data_source_0/data_index[0]_net_1 ), .B(
        \data_source_0/data_index[8]_net_1 ), .C(
        \data_source_0/tag_control_sig_2_0_a20_0[7] ), .Y(
        \data_source_0/N_927 ));
    NOR2B \switching_circuit_0/un180_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[18] ), .B(
        main_clock_0_clock_out), .Y(
        \switching_circuit_0/un180_out_signal_switch_0_net_1 ));
    NOR2B \data_source_0/data_index_RNIBM6D[4]  (.A(
        \data_source_0/N_668 ), .B(\data_source_0/data_index[4]_net_1 )
        , .Y(\data_source_0/N_901_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_7[4]  (.D(
        \data_source_0/tag_data_buf_7_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_7[4]_net_1 ));
    AND3 \data_source_0/un3_data_index_I_24  (.A(
        \data_source_0/DWACT_FINC_E[0] ), .B(
        \data_source_0/DWACT_FINC_E[2] ), .C(
        \data_source_0/DWACT_FINC_E[3] ), .Y(
        \data_source_0/DWACT_FINC_E[4] ));
    NOR2B \data_source_0/data_index_RNIRO0M[7]  (.A(
        \data_source_0/N_1143 ), .B(\data_source_0/N_1141 ), .Y(
        \data_source_0/N_1163 ));
    AO1 \data_source_0/data_index_RNINCII2[2]  (.A(
        \data_source_0/N_1189 ), .B(\data_source_0/N_1181 ), .C(
        \data_source_0/N_1221 ), .Y(\data_source_0/N_764 ));
    NOR2B \data_source_0/tag_data_buf_12_RNO[6]  (.A(
        \data_source_0/tag_data_buf_12[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_12_4[6] ));
    AND3 \main_clock_0/un5_counter_1_I_18  (.A(
        \main_clock_0/counter[3]_net_1 ), .B(
        \main_clock_0/counter[4]_net_1 ), .C(
        \main_clock_0/counter[5]_net_1 ), .Y(
        \main_clock_0/DWACT_FINC_E[2] ));
    NOR2B \data_source_0/tag_data_buf_16_RNIF69P[7]  (.A(
        \data_source_0/tag_data_buf_16[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[15] ));
    XA1A \switching_circuit_0/un13_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[1] ), 
        .C(\data_source_0_tag_control_sig[1] ), .Y(
        \switching_circuit_0/un13_out_signal_switch_0_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_5[8]  (.A(
        \data_source_0/N_1210 ), .B(\data_source_0/N_1181 ), .Y(
        \data_source_0/N_955 ));
    XOR2 \main_clock_0/un5_counter_1_I_20  (.A(\main_clock_0/N_2 ), .B(
        \main_clock_0/counter[7]_net_1 ), .Y(\main_clock_0/I_20_0 ));
    OA1 \data_source_0/tag_control_sig_RNO_16[18]  (.A(
        \data_source_0/N_1227 ), .B(\data_source_0/N_1232 ), .C(
        \data_source_0/N_1186 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_1_0[18] ));
    CLKINT \main_clock_0/clock_out_RNIG44  (.A(
        \main_clock_0/clock_out_i ), .Y(main_clock_0_clock_out));
    DFN1C0 \main_clock_0/counter[4]  (.D(\main_clock_0/I_12_0 ), .CLK(
        GLA), .CLR(reset_c), .Q(\main_clock_0/counter[4]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_16_RNO[1]  (.A(
        \data_source_0/tag_data_buf_16[0]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_16_4[1] ));
    NOR2B \data_source_0/data_index_RNID81C1_0[5]  (.A(
        \data_source_0/N_1183 ), .B(\data_source_0/N_1161 ), .Y(
        \data_source_0/N_835 ));
    NOR2B \data_source_0/data_index_RNIIMJH_2[0]  (.A(
        \data_source_0/N_1144 ), .B(\data_source_0/N_1132 ), .Y(
        \data_source_0/N_1173 ));
    NOR3B \data_source_0/tag_control_sig_RNO_14[6]  (.A(
        \data_source_0/N_1144 ), .B(
        \data_source_0/tag_control_sig_2_0_a20_2_0[6] ), .C(
        \data_source_0/data_index[3]_net_1 ), .Y(\data_source_0/N_917 )
        );
    NOR2B \data_source_0/data_index_0_RNIJ6UA1[7]  (.A(
        \data_source_0/N_1198 ), .B(\data_source_0/N_1190 ), .Y(
        \data_source_0/N_1218 ));
    AO1 \data_source_0/tag_control_sig_RNO_4[9]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_2_0[9] ), .B(
        \data_source_0/N_1239 ), .C(\data_source_0/N_964 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[9] ));
    NOR2B \data_source_0/tag_control_sig_RNO_21[1]  (.A(
        \data_source_0/N_1199 ), .B(\data_source_0/N_1186 ), .Y(
        \data_source_0/N_847 ));
    AO1 \data_source_0/tag_control_sig_RNO_9[5]  (.A(
        \data_source_0/N_1192 ), .B(\data_source_0/N_1186 ), .C(
        \data_source_0/N_904 ), .Y(
        \data_source_0/tag_control_sig_2_0_4[5] ));
    NOR2B \data_source_0/tag_data_buf_15_RNO[7]  (.A(
        \data_source_0/tag_data_buf_15[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_15_4[7] ));
    DFN1E1C0 \data_source_0/tag_data_buf_15[7]  (.D(
        \data_source_0/tag_data_buf_15_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_15[7]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_11[7]  (.D(
        \data_source_0/tag_data_buf_11_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_11[7]_net_1 ));
    OR2 \modulator_0/output_signal_RNO_7  (.A(
        \modulator_0/clock_counter[5]_net_1 ), .B(
        \modulator_0/clock_counter[4]_net_1 ), .Y(
        \modulator_0/un5lto5 ));
    NOR2B \data_source_0/tag_control_sig_RNO_4[2]  (.A(
        \data_source_0/N_1226 ), .B(\data_source_0/N_1177 ), .Y(
        \data_source_0/N_859 ));
    AX1C \data_source_0/un3_data_index_I_26  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/DWACT_FINC_E[4] ), .C(
        \data_source_0/data_index[9]_net_1 ), .Y(\data_source_0/I_26 ));
    AO1 \data_source_0/tag_control_sig_RNO_9[13]  (.A(
        \data_source_0/N_1196 ), .B(\data_source_0/N_1177 ), .C(
        \data_source_0/N_1031 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[13] ));
    NOR2A \data_source_0/data_index_RNI3LP8_1[0]  (.A(
        \data_source_0/data_index[3]_net_1 ), .B(
        \data_source_0/data_index[0]_net_1 ), .Y(
        \data_source_0/N_1142 ));
    XOR2 \data_source_0/un3_data_index_I_14  (.A(\data_source_0/N_6 ), 
        .B(\data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/I_14 ));
    NOR2A \data_source_0/data_index_RNI3LP8_2[0]  (.A(
        \data_source_0/data_index[0]_net_1 ), .B(
        \data_source_0/data_index[3]_net_1 ), .Y(
        \data_source_0/N_1132 ));
    DFN1E1C0 \data_source_0/tag_data_buf_11[2]  (.D(
        \data_source_0/tag_data_buf_11_4[2] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_11[2]_net_1 ));
    XOR2 \data_source_0/data_index_RNI6OP8[0]  (.A(
        \data_source_0/data_index[0]_net_1 ), .B(
        \data_source_0/data_index[6]_net_1 ), .Y(
        \data_source_0/N_703_i ));
    NOR2B \data_source_0/tag_control_sig_RNO_19[14]  (.A(
        \data_source_0/N_1202 ), .B(\data_source_0/N_1179 ), .Y(
        \data_source_0/N_1049 ));
    DFN1E1C0 \data_source_0/tag_data_buf_1[4]  (.D(
        \data_source_0/tag_data_buf_1_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_1[4]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_21[5]  (.A(
        \data_source_0/N_1173 ), .B(\data_source_0/N_1180 ), .C(
        \data_source_0/N_1160 ), .Y(\data_source_0/N_807 ));
    OA1 \data_source_0/tag_control_sig_RNO_19[1]  (.A(
        \data_source_0/N_1179 ), .B(\data_source_0/N_1178 ), .C(
        \data_source_0/N_1216 ), .Y(\data_source_0/N_829 ));
    NOR2B \switching_circuit_0/un80_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[8] ), .B(main_clock_0_clock_out)
        , .Y(\switching_circuit_0/un80_out_signal_switch_0_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_5[13]  (.A(
        \data_source_0/N_1035 ), .B(\data_source_0/N_1025 ), .C(
        \data_source_0/tag_control_sig_2_0_1[13] ), .Y(
        \data_source_0/tag_control_sig_2_0_10[13] ));
    DFN1E1C0 \modulator_0/clock_counter[9]  (.D(
        \modulator_0/clock_counter_n9 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/un6lto9 ));
    DFN1E1C0 \data_source_0/tag_data_buf_7[7]  (.D(
        \data_source_0/tag_data_buf_7_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_7[7]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_3_RNO[3]  (.A(
        \data_source_0/tag_data_buf_3[2]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_3_4[3] ));
    NOR2B \data_source_0/tag_data_buf_1_RNO[6]  (.A(
        \data_source_0/tag_data_buf_1[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_1_4[6] ));
    OR2 \data_source_0/tag_control_sig_RNO_11[8]  (.A(
        \data_source_0/N_1193 ), .B(\data_source_0/N_1180 ), .Y(
        \data_source_0/N_800 ));
    DFN1E1 \data_source_0/tag_control_sig[5]  (.D(
        \data_source_0/tag_control_sig_2[5] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[5] ));
    OR3 \data_source_0/tag_control_sig_RNO_2[9]  (.A(
        \data_source_0/tag_control_sig_2_0_3[9] ), .B(
        \data_source_0/tag_control_sig_2_0_2[9] ), .C(
        \data_source_0/tag_control_sig_2_0_11[9] ), .Y(
        \data_source_0/tag_control_sig_2_0_14[9] ));
    NOR2B \data_source_0/tag_control_sig_RNO_4[15]  (.A(
        \data_source_0/N_1213 ), .B(\data_source_0/N_1199 ), .Y(
        \data_source_0/N_1062 ));
    NOR2B \data_source_0/tag_control_sig_RNO_15[19]  (.A(
        \data_source_0/N_1199 ), .B(\data_source_0/N_1185 ), .Y(
        \data_source_0/N_1125 ));
    AO1 \data_source_0/tag_control_sig_RNO_7[19]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_0_0[19] ), .B(
        \data_source_0/N_1074_2 ), .C(\data_source_0/N_1129 ), .Y(
        \data_source_0/tag_control_sig_2_0_2[19] ));
    DFN1E1 \data_source_0/tag_control_sig[18]  (.D(
        \data_source_0/tag_control_sig_2[18] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[18] ));
    IOPAD_TRI \output_signal_pad[3]/U0/U0  (.D(
        \output_signal_pad[3]/U0/NET1 ), .E(
        \output_signal_pad[3]/U0/NET2 ), .PAD(output_signal[3]));
    NOR2B \data_source_0/tag_control_sig_RNO_18[11]  (.A(
        \data_source_0/N_1226 ), .B(\data_source_0/N_1160 ), .Y(
        \data_source_0/N_990 ));
    NOR2 \data_source_0/data_index_RNI8J6D[1]  (.A(
        \data_source_0/N_668 ), .B(\data_source_0/data_index[1]_net_1 )
        , .Y(\data_source_0/N_1040_1 ));
    NOR2B \data_source_0/data_index_RNI46K71[6]  (.A(
        \data_source_0/N_1195 ), .B(\data_source_0/N_1178 ), .Y(
        \data_source_0/N_1027 ));
    AO1 \data_source_0/tag_control_sig_2_0_4[15]  (.A(
        \data_source_0/N_1175 ), .B(\data_source_0/N_1206 ), .C(
        \data_source_0/N_1042 ), .Y(
        \data_source_0/tag_control_sig_2_0_4[15]_net_1 ));
    XA1A \data_source_0/counter_RNO[11]  (.A(\data_source_0/N_40 ), .B(
        \data_source_0/counter[11]_net_1 ), .C(
        modulator_0_output_signal), .Y(\data_source_0/counter_n11 ));
    NOR2B \modulator_0/clock_counter_RNI3U8B[8]  (.A(
        \modulator_0/clock_counter_c7 ), .B(
        \modulator_0/clock_counter[8]_net_1 ), .Y(
        \modulator_0/clock_counter_c8 ));
    NOR2B \data_source_0/tag_data_buf_17_RNO[1]  (.A(
        \data_source_0/tag_data_buf_17[0]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_17_4[1] ));
    NOR2B \switching_circuit_0/un120_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[12] ), .B(
        main_clock_0_clock_out), .Y(
        \switching_circuit_0/un120_out_signal_switch_0_net_1 ));
    AOI1B \data_source_0/data_index_RNO[1]  (.A(
        \data_source_0/tag_control_sig_1_649_6 ), .B(
        \data_source_0/tag_control_sig_1_3[649] ), .C(
        \data_source_0/I_5 ), .Y(\data_source_0/data_index_3[1] ));
    NOR2B \data_source_0/tag_data_buf_19_RNO[5]  (.A(
        \data_source_0/tag_data_buf_19[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_19_4[5] ));
    NOR2B \data_source_0/data_index_RNIIF0M_9[6]  (.A(
        \data_source_0/N_1148 ), .B(\data_source_0/N_1140 ), .Y(
        \data_source_0/N_1196 ));
    DFN1E1C0 \data_source_0/tag_data_buf_11[6]  (.D(
        \data_source_0/tag_data_buf_11_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_11[6]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_7[6]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_1_0[6] ), .B(
        \data_source_0/N_1179 ), .C(\data_source_0/N_917 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[6] ));
    NOR2B \data_source_0/tag_control_sig_RNO_19[9]  (.A(
        \data_source_0/N_1195 ), .B(\data_source_0/N_1181 ), .Y(
        \data_source_0/N_968 ));
    NOR3B \data_source_0/tag_control_sig_RNO_18[6]  (.A(
        \data_source_0/N_1148 ), .B(\data_source_0/N_704_i ), .C(
        \data_source_0/data_index_0[4]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_2_0[6] ));
    NOR3C \data_source_0/tag_control_sig_RNO_12[16]  (.A(
        \data_source_0/N_759 ), .B(\data_source_0/N_1142 ), .C(
        \data_source_0/tag_control_sig_2_0_a20_2[16] ), .Y(
        \data_source_0/N_1072 ));
    NOR2B \switching_circuit_0/un100_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[10] ), .B(
        main_clock_0_clock_out), .Y(
        \switching_circuit_0/un100_out_signal_switch_0_net_1 ));
    AND3 \data_source_0/un3_data_index_I_16  (.A(
        \data_source_0/DWACT_FINC_E[0] ), .B(
        \data_source_0/DWACT_FINC_E[1] ), .C(
        \data_source_0/data_index[5]_net_1 ), .Y(\data_source_0/N_5 ));
    OR2A \data_source_0/tag_data_buf_2_RNO[1]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_2[0]_net_1 ), .Y(
        \data_source_0/tag_data_buf_2_4[1] ));
    OR2A \data_source_0/tag_data_buf_6_RNO[1]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_6[0]_net_1 ), .Y(
        \data_source_0/tag_data_buf_6_4[1] ));
    NOR3C \data_source_0/tag_control_sig_RNO_20[17]  (.A(
        \data_source_0/N_1140 ), .B(\data_source_0/N_1154 ), .C(
        \data_source_0/N_1179 ), .Y(\data_source_0/N_1097 ));
    XA1A \data_source_0/counter_RNO[12]  (.A(\data_source_0/N_41 ), .B(
        \data_source_0/counter[12]_net_1 ), .C(
        modulator_0_output_signal), .Y(\data_source_0/counter_n12 ));
    NOR2B \data_source_0/tag_data_buf_14_RNO[7]  (.A(
        \data_source_0/tag_data_buf_14[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_14_4[7] ));
    NOR3C \data_source_0/tag_control_sig_RNO_7[12]  (.A(
        \data_source_0/N_1156 ), .B(\data_source_0/N_1155 ), .C(
        \data_source_0/N_1177 ), .Y(\data_source_0/N_1019 ));
    OR3 \data_source_0/tag_control_sig_RNO_11[14]  (.A(
        \data_source_0/N_1040 ), .B(\data_source_0/N_1049 ), .C(
        \data_source_0/tag_control_sig_2_0_3[14] ), .Y(
        \data_source_0/tag_control_sig_2_0_10[14] ));
    AO1 \data_source_0/tag_control_sig_RNO_15[15]  (.A(
        \data_source_0/N_1209 ), .B(\data_source_0/N_1181 ), .C(
        \data_source_0/N_1066 ), .Y(
        \data_source_0/tag_control_sig_2_0_2[15] ));
    OR3 \data_source_0/tag_control_sig_RNO[16]  (.A(
        \data_source_0/tag_control_sig_2_0_9[16] ), .B(
        \data_source_0/tag_control_sig_2_0_8[16] ), .C(
        \data_source_0/tag_control_sig_2_0_13[16] ), .Y(
        \data_source_0/tag_control_sig_2[16] ));
    AO1 \data_source_0/tag_control_sig_RNO_20[13]  (.A(
        \data_source_0/N_1200 ), .B(\data_source_0/N_1163 ), .C(
        \data_source_0/N_1034 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[13] ));
    DFN1E1C0 \data_source_0/tag_data_buf_10[7]  (.D(
        \data_source_0/tag_data_buf_10_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_10[7]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_21[7]  (.A(
        \data_source_0/N_1156 ), .B(
        \data_source_0/data_index[9]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_4_1[7] ));
    OR2 \data_source_0/tag_control_sig_RNO[7]  (.A(
        \data_source_0/tag_control_sig_2_0_12[7] ), .B(
        \data_source_0/tag_control_sig_2_0_11[7] ), .Y(
        \data_source_0/tag_control_sig_2[7] ));
    DFN1E1C0 \data_source_0/tag_data_buf_5[5]  (.D(
        \data_source_0/tag_data_buf_5_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_5[5]_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_18[8]  (.A(
        \data_source_0/N_1142 ), .B(
        \data_source_0/data_index[7]_net_1 ), .C(
        \data_source_0/N_1211 ), .Y(\data_source_0/N_950 ));
    DFN1E1P0 \data_source_0/tag_data_buf_19[1]  (.D(
        \data_source_0/tag_data_buf_19_4[1] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_19[1]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_17_RNO[6]  (.A(
        \data_source_0/tag_data_buf_17[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_17_4[6] ));
    OR2 \data_source_0/tag_control_sig_RNO_6[10]  (.A(
        \data_source_0/N_755 ), .B(\data_source_0/N_1162 ), .Y(
        \data_source_0/N_779 ));
    OR3 \data_source_0/tag_control_sig_RNO_0[8]  (.A(
        \data_source_0/N_945 ), .B(\data_source_0/N_879 ), .C(
        \data_source_0/tag_control_sig_2_0_3[8] ), .Y(
        \data_source_0/tag_control_sig_2_0_9[8] ));
    NOR2B \data_source_0/tag_data_buf_16_RNO[7]  (.A(
        \data_source_0/tag_data_buf_16[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_16_4[7] ));
    NOR2A \modulator_0/counter_RNO[0]  (.A(
        \modulator_0/counter_0_sqmuxa ), .B(
        \modulator_0/counter[0]_net_1 ), .Y(\modulator_0/counter_n0 ));
    DFN1E1C0 \data_source_0/tag_data_buf_18[5]  (.D(
        \data_source_0/tag_data_buf_18_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_18[5]_net_1 ));
    NOR2B \data_source_0/data_index_RNI46K71_0[6]  (.A(
        \data_source_0/N_1201 ), .B(\data_source_0/N_1184 ), .Y(
        \data_source_0/N_819 ));
    DFN1C0 \modulator_0/counter[5]  (.D(\modulator_0/counter_n5 ), 
        .CLK(main_clock_0_clock_out), .CLR(reset_c), .Q(
        \modulator_0/counter[5]_net_1 ));
    XOR2 \data_source_0/un3_data_index_I_23  (.A(\data_source_0/N_3 ), 
        .B(\data_source_0/data_index[8]_net_1 ), .Y(
        \data_source_0/I_23 ));
    NOR2 \data_source_0/data_index_RNIASP8_0[4]  (.A(
        \data_source_0/data_index[6]_net_1 ), .B(
        \data_source_0/data_index[4]_net_1 ), .Y(
        \data_source_0/N_1135 ));
    NOR2B \switching_circuit_0/un60_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[6] ), .B(main_clock_0_clock_out)
        , .Y(\switching_circuit_0/un60_out_signal_switch_0_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_18[2]  (.D(
        \data_source_0/tag_data_buf_18_4[2] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_18[2]_net_1 ));
    XOR2 \data_source_0/un3_data_index_I_9  (.A(\data_source_0/N_8 ), 
        .B(\data_source_0/data_index[3]_net_1 ), .Y(
        \data_source_0/I_9 ));
    DFN1E1C0 \data_source_0/tag_data_buf_2[6]  (.D(
        \data_source_0/tag_data_buf_2_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_2[6]_net_1 ));
    MX2 \switching_circuit_0/out_signal_switch_1[4]  (.A(
        \switching_circuit_0/un40_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un43_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[4] ));
    AO1 \data_source_0/tag_control_sig_RNO_15[13]  (.A(
        \data_source_0/N_1192 ), .B(\data_source_0/N_1182 ), .C(
        \data_source_0/N_1021 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[13] ));
    NOR3C \data_source_0/data_index_RNIJ6UA1[6]  (.A(
        \data_source_0/tag_control_sig_1_3[649] ), .B(
        \data_source_0/N_1148 ), .C(\data_source_0/N_1179 ), .Y(
        \data_source_0/N_1220 ));
    NOR2B \switching_circuit_0/un160_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[16] ), .B(
        main_clock_0_clock_out), .Y(
        \switching_circuit_0/un160_out_signal_switch_0_net_1 ));
    XA1A \switching_circuit_0/un113_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[11] ), 
        .C(\data_source_0_tag_control_sig[11] ), .Y(
        \switching_circuit_0/un113_out_signal_switch_0_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO[4]  (.A(
        \data_source_0/tag_control_sig_2_0_9[4] ), .B(
        \data_source_0/tag_control_sig_2_0_8[4] ), .C(
        \data_source_0/tag_control_sig_2_0_13[4] ), .Y(
        \data_source_0/tag_control_sig_2[4] ));
    NOR2A \data_source_0/data_index_RNIB80M[3]  (.A(
        \data_source_0/N_1238 ), .B(\data_source_0/N_704_i ), .Y(
        \data_source_0/N_1074_2 ));
    AO1 \data_source_0/tag_control_sig_RNO_17[19]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_12_0[19] ), .B(
        \data_source_0/N_1237 ), .C(\data_source_0/N_1122 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[19] ));
    OR3 \data_source_0/tag_control_sig_RNO_0[15]  (.A(
        \data_source_0/tag_control_sig_2_0_0[15] ), .B(
        \data_source_0/N_1062 ), .C(
        \data_source_0/tag_control_sig_2_0_10[15] ), .Y(
        \data_source_0/tag_control_sig_2_0_14[15] ));
    DFN1E1C0 \data_source_0/tag_data_buf_14[4]  (.D(
        \data_source_0/tag_data_buf_14_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_14[4]_net_1 ));
    NOR2B \data_source_0/data_index_RNIFQ6D[5]  (.A(
        \data_source_0/N_1135 ), .B(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/N_1151 ));
    IOPAD_TRI \output_signal_pad[17]/U0/U0  (.D(
        \output_signal_pad[17]/U0/NET1 ), .E(
        \output_signal_pad[17]/U0/NET2 ), .PAD(output_signal[17]));
    AO1 \data_source_0/tag_control_sig_RNO_9[8]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_6_0[7] ), .B(
        \data_source_0/N_1191 ), .C(\data_source_0/N_947 ), .Y(
        \data_source_0/tag_control_sig_2_0_4[8] ));
    NOR3B \data_source_0/tag_control_sig_RNO_12[17]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/data_index[3]_net_1 ), .C(
        \data_source_0/data_index_0[7]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_2_1[17] ));
    AOI1D \data_source_0/tag_control_sig_RNO_19[18]  (.A(
        \data_source_0/N_1162 ), .B(\data_source_0/N_1159 ), .C(
        \data_source_0/N_1190 ), .Y(\data_source_0/N_1102 ));
    NOR3B \data_source_0/tag_control_sig_RNO_16[16]  (.A(
        \data_source_0/N_1182 ), .B(\data_source_0/N_1183 ), .C(
        \data_source_0/data_index_0[7]_net_1 ), .Y(
        \data_source_0/N_1081 ));
    NOR3C \data_source_0/data_index_RNIJ6UA1_0[2]  (.A(
        \data_source_0/N_1156 ), .B(\data_source_0/N_1155 ), .C(
        \data_source_0/N_1185 ), .Y(\data_source_0/N_1221 ));
    NOR2B \data_source_0/tag_control_sig_RNO_13[17]  (.A(
        \data_source_0/N_1145 ), .B(\data_source_0/N_1192 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_0_0[17] ));
    NOR2B \data_source_0/data_index_RNI1V0M[7]  (.A(
        \data_source_0/N_1143 ), .B(\data_source_0/N_1134 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_3_0[9] ));
    DFN1E1P0 \data_source_0/tag_data_buf_5[0]  (.D(
        \data_source_0/tag_data_buf_5_4[0] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_5[0]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_7_RNO[5]  (.A(
        \data_source_0/tag_data_buf_7[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_7_4[5] ));
    OR3 \data_source_0/tag_control_sig_RNO[17]  (.A(
        \data_source_0/tag_control_sig_2_0_10[17] ), .B(
        \data_source_0/tag_control_sig_2_0_9[17] ), .C(
        \data_source_0/tag_control_sig_2_0_14[17] ), .Y(
        \data_source_0/tag_control_sig_2[17] ));
    AND2 \data_source_0/tag_control_sig_2_0_a20_13[11]  (.A(
        \data_source_0/N_1181 ), .B(\data_source_0/N_1200 ), .Y(
        \data_source_0/N_1001 ));
    OR3 \data_source_0/tag_control_sig_RNO_2[6]  (.A(
        \data_source_0/tag_control_sig_2_0_9[6] ), .B(
        \data_source_0/tag_control_sig_2_0_8[6] ), .C(
        \data_source_0/tag_control_sig_2_0_12[6] ), .Y(
        \data_source_0/tag_control_sig_2_0_15[6] ));
    NOR2B \data_source_0/data_index_RNIIF0M[4]  (.A(
        \data_source_0/N_1148 ), .B(\data_source_0/N_1134 ), .Y(
        \data_source_0/N_1190 ));
    AO1 \data_source_0/tag_control_sig_RNO_4[4]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_8_0[4] ), .B(
        \data_source_0/N_1163 ), .C(
        \data_source_0/tag_control_sig_RNO_11[4]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[4] ));
    AO1 \data_source_0/tag_control_sig_RNO_3[2]  (.A(
        \data_source_0/N_1225 ), .B(\data_source_0/N_1176 ), .C(
        \data_source_0/N_860 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[2] ));
    XA1A \switching_circuit_0/un93_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[9] ), 
        .C(\data_source_0_tag_control_sig[9] ), .Y(
        \switching_circuit_0/un93_out_signal_switch_0_net_1 ));
    NOR3B \data_source_0/tag_control_sig_RNO_17[15]  (.A(
        \data_source_0/N_1182 ), .B(
        \data_source_0/tag_control_sig_2_0_a20_0_1[15] ), .C(
        \data_source_0/N_707_i ), .Y(\data_source_0/N_1055 ));
    NOR3C \data_source_0/tag_control_sig_RNO_13[3]  (.A(
        \data_source_0/N_1140 ), .B(\data_source_0/N_1154 ), .C(
        \data_source_0/N_780 ), .Y(\data_source_0/N_865 ));
    NOR2B \data_source_0/data_index_RNI3LP8_0[0]  (.A(
        \data_source_0/data_index[0]_net_1 ), .B(
        \data_source_0/data_index[3]_net_1 ), .Y(
        \data_source_0/N_1138 ));
    XA1A \switching_circuit_0/un53_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[5] ), 
        .C(\data_source_0_tag_control_sig[5] ), .Y(
        \switching_circuit_0/un53_out_signal_switch_0_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_7[16]  (.A(
        \data_source_0/N_1208 ), .B(\data_source_0/N_1163 ), .C(
        \data_source_0/N_1040_1 ), .Y(\data_source_0/N_1076 ));
    NOR3B \data_source_0/tag_control_sig_RNO_15[9]  (.A(
        \data_source_0/N_1149 ), .B(\data_source_0/N_919_1 ), .C(
        \data_source_0/data_index_0[4]_net_1 ), .Y(
        \data_source_0/N_961 ));
    IOPAD_IN \mac_control_signal_pad/U0/U0  (.PAD(mac_control_signal), 
        .Y(\mac_control_signal_pad/U0/NET1 ));
    NOR3C \modulator_0/counter_RNINTKF1[2]  (.A(
        \modulator_0/counter[1]_net_1 ), .B(
        \modulator_0/counter[0]_net_1 ), .C(
        \modulator_0/counter[2]_net_1 ), .Y(\modulator_0/counter_c2 ));
    AND3 \data_source_0/un3_data_index_I_13  (.A(
        \data_source_0/DWACT_FINC_E[0] ), .B(
        \data_source_0/data_index[3]_net_1 ), .C(
        \data_source_0/data_index_0[4]_net_1 ), .Y(\data_source_0/N_6 )
        );
    AOI1B \data_source_0/data_index_RNO[9]  (.A(
        \data_source_0/tag_control_sig_1_649_6 ), .B(
        \data_source_0/tag_control_sig_1_3[649] ), .C(
        \data_source_0/I_26 ), .Y(\data_source_0/data_index_3[9] ));
    NOR2B \data_source_0/data_index_RNIIF0M_7[6]  (.A(
        \data_source_0/tag_control_sig_1_3[649] ), .B(
        \data_source_0/N_1154 ), .Y(\data_source_0/N_1209 ));
    NOR2B \data_source_0/tag_control_sig_RNO_7[11]  (.A(
        \data_source_0/N_1206 ), .B(\data_source_0/N_1163 ), .Y(
        \data_source_0/N_991 ));
    OR2A \data_source_0/tag_data_buf_3_RNO[0]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_3[7]_net_1 ), .Y(
        \data_source_0/tag_data_buf_3_4[0] ));
    DFN1C0 \data_source_0/counter[8]  (.D(\data_source_0/N_12 ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .Q(
        \data_source_0/counter[8]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_6[0]  (.D(
        \data_source_0/output_data_23[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_6[0]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_0[7]  (.A(
        \data_source_0/tag_control_sig_2_0_6[7] ), .B(
        \data_source_0/tag_control_sig_2_0_5[7] ), .C(
        \data_source_0/tag_control_sig_2_0_9[7] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[7] ));
    DFN1E1C0 \data_source_0/tag_data_buf_1[5]  (.D(
        \data_source_0/tag_data_buf_1_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_1[5]_net_1 ));
    OA1 \data_source_0/tag_control_sig_RNO_6[4]  (.A(
        \data_source_0/N_783 ), .B(\data_source_0/N_996_1 ), .C(
        \data_source_0/N_1204 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[4] ));
    NOR2B \switching_circuit_0/un1_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[0] ), .B(main_clock_0_clock_out)
        , .Y(\switching_circuit_0/un1_out_signal_switch_0_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_21[8]  (.A(
        \data_source_0/N_1152 ), .B(\data_source_0/N_1175 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_6_0[8] ));
    NOR3B \data_source_0/tag_control_sig_RNO_6[17]  (.A(
        \data_source_0/N_1180 ), .B(
        \data_source_0/tag_control_sig_2_0_a20_4_1[17] ), .C(
        \data_source_0/N_701_i ), .Y(\data_source_0/N_1091 ));
    DFN1E1C0 \data_source_0/output_data[13]  (.D(
        \data_source_0/output_data_23[13] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[13] ));
    NOR2 \main_clock_0/counter_RNIF4VS[1]  (.A(
        \main_clock_0/counter[4]_net_1 ), .B(
        \main_clock_0/counter[1]_net_1 ), .Y(
        \main_clock_0/counter14_2 ));
    OR2A \data_source_0/tag_data_buf_13_RNO[3]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_13[2]_net_1 ), .Y(
        \data_source_0/tag_data_buf_13_4[3] ));
    NOR2A \data_source_0/tag_control_sig_RNO_11[18]  (.A(
        \data_source_0/N_1155 ), .B(
        \data_source_0/data_index[4]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_2_0[18] ));
    AO1 \modulator_0/output_signal_RNO_1  (.A(\modulator_0/un6lt11 ), 
        .B(\modulator_0/un6lto11 ), .C(\modulator_0/un6lto12 ), .Y(
        \modulator_0/un6lt15 ));
    NOR2B \data_source_0/tag_data_buf_8_RNO[4]  (.A(
        \data_source_0/tag_data_buf_8[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_8_4[4] ));
    NOR3C \data_source_0/tag_control_sig_RNO_17[13]  (.A(
        \data_source_0/N_1140 ), .B(\data_source_0/N_1154 ), .C(
        \data_source_0/N_1173 ), .Y(\data_source_0/N_1031 ));
    NOR2B \data_source_0/tag_data_buf_19_RNO[6]  (.A(
        \data_source_0/tag_data_buf_19[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_19_4[6] ));
    DFN1E1C0 \data_source_0/tag_data_buf_18[7]  (.D(
        \data_source_0/tag_data_buf_18_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_18[7]_net_1 ));
    OR2A \data_source_0/tag_data_buf_19_RNO[0]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_19[7]_net_1 ), .Y(
        \data_source_0/tag_data_buf_19_4[0] ));
    AO1 \data_source_0/tag_control_sig_RNO_20[14]  (.A(
        \data_source_0/N_1206 ), .B(\data_source_0/N_1180 ), .C(
        \data_source_0/N_1045 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[14] ));
    IOTRI_OB_EB \output_signal_pad[11]/U0/U1  (.D(
        \output_signal_c[11] ), .E(VCC), .DOUT(
        \output_signal_pad[11]/U0/NET1 ), .EOUT(
        \output_signal_pad[11]/U0/NET2 ));
    IOPAD_TRI \output_signal_pad[18]/U0/U0  (.D(
        \output_signal_pad[18]/U0/NET1 ), .E(
        \output_signal_pad[18]/U0/NET2 ), .PAD(output_signal[18]));
    OR2A \data_source_0/tag_data_buf_13_RNO[2]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_13[1]_net_1 ), .Y(
        \data_source_0/tag_data_buf_13_4[2] ));
    XA1A \switching_circuit_0/un153_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[15] ), 
        .C(\data_source_0_tag_control_sig[15] ), .Y(
        \switching_circuit_0/un153_out_signal_switch_0_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_18[12]  (.A(
        \data_source_0/N_707_i ), .B(\data_source_0/N_1161 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_1_0[12] ));
    NOR3C \data_source_0/tag_control_sig_RNO_16[17]  (.A(
        \data_source_0/N_1178 ), .B(\data_source_0/N_668 ), .C(
        \data_source_0/N_1227 ), .Y(\data_source_0/N_1092 ));
    NOR3A \data_source_0/tag_control_sig_RNO_13[5]  (.A(
        \data_source_0/N_1148 ), .B(
        \data_source_0/data_index_0[4]_net_1 ), .C(
        \data_source_0/N_704_i ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_1_0[5] ));
    IOTRI_OB_EB \signal_into_switch_pad/U0/U1  (.D(VCC), .E(VCC), 
        .DOUT(\signal_into_switch_pad/U0/NET1 ), .EOUT(
        \signal_into_switch_pad/U0/NET2 ));
    AO1 \data_source_0/tag_control_sig_RNO_9[15]  (.A(
        \data_source_0/N_1201 ), .B(\data_source_0/N_1180 ), .C(
        \data_source_0/N_1055 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[15] ));
    IOPAD_TRI \output_signal_pad[10]/U0/U0  (.D(
        \output_signal_pad[10]/U0/NET1 ), .E(
        \output_signal_pad[10]/U0/NET2 ), .PAD(output_signal[10]));
    DFN1E1C0 \data_source_0/tag_data_buf_13[6]  (.D(
        \data_source_0/tag_data_buf_13_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_13[6]_net_1 ));
    DFN1E1P0 \data_source_0/tag_data_buf_10[1]  (.D(
        \data_source_0/tag_data_buf_10_4[1] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_10[1]_net_1 ));
    OR2A \data_source_0/data_index_0_RNIQT3C[4]  (.A(
        \data_source_0/data_index[7]_net_1 ), .B(
        \data_source_0/data_index_0[4]_net_1 ), .Y(
        \data_source_0/N_759 ));
    IOPAD_TRI \output_signal_pad[13]/U0/U0  (.D(
        \output_signal_pad[13]/U0/NET1 ), .E(
        \output_signal_pad[13]/U0/NET2 ), .PAD(output_signal[13]));
    NOR2B \data_source_0/output_data_RNO[10]  (.A(
        \data_source_0/tag_data_buf_11[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[10] ));
    DFN1C0 \main_clock_0/counter[7]  (.D(\main_clock_0/I_20_0 ), .CLK(
        GLA), .CLR(reset_c), .Q(\main_clock_0/counter[7]_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_15[10]  (.A(
        \data_source_0/N_1133 ), .B(\data_source_0/N_1151 ), .C(
        \data_source_0/N_1198 ), .Y(\data_source_0/N_982 ));
    OR3 \data_source_0/tag_control_sig_RNO_1[4]  (.A(
        \data_source_0/N_881 ), .B(\data_source_0/N_764 ), .C(
        \data_source_0/tag_control_sig_2_0_0[4] ), .Y(
        \data_source_0/tag_control_sig_2_0_8[4] ));
    DFN1E1C0 \data_source_0/tag_data_buf_6[7]  (.D(
        \data_source_0/tag_data_buf_6_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_6[7]_net_1 ));
    NOR2B \data_source_0/data_index_RNIIF0M_1[6]  (.A(
        \data_source_0/N_1147 ), .B(\data_source_0/N_1136 ), .Y(
        \data_source_0/N_1195 ));
    DFN1E1C0 \data_source_0/tag_data_buf_12[5]  (.D(
        \data_source_0/tag_data_buf_12_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_12[5]_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_13[0]  (.A(
        \data_source_0/N_1173 ), .B(
        \data_source_0/tag_control_sig_1_3[649] ), .C(
        \data_source_0/N_1233 ), .Y(\data_source_0/N_815 ));
    INV \data_source_0/un3_data_index_I_4  (.A(
        \data_source_0/data_index[0]_net_1 ), .Y(\data_source_0/I_4 ));
    MX2 \switching_circuit_0/out_signal_switch_1[15]  (.A(
        \switching_circuit_0/un150_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un153_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[15] ));
    OR3 \data_source_0/tag_control_sig_RNO_5[15]  (.A(
        \data_source_0/N_1068 ), .B(\data_source_0/N_1057 ), .C(
        \data_source_0/tag_control_sig_2_0_2[15] ), .Y(
        \data_source_0/tag_control_sig_2_0_10[15] ));
    NOR2B \data_source_0/tag_data_buf_7_RNO[4]  (.A(
        \data_source_0/tag_data_buf_7[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_7_4[4] ));
    DFN1E1C0 \data_source_0/tag_data_buf_8[2]  (.D(
        \data_source_0/tag_data_buf_8_4[2] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_8[2]_net_1 ));
    NOR2A \data_source_0/data_index_RNI3LP8_1[1]  (.A(
        \data_source_0/data_index[2]_net_1 ), .B(
        \data_source_0/data_index[1]_net_1 ), .Y(
        \data_source_0/N_1152 ));
    AOI1B \modulator_0/output_signal_RNO  (.A(\modulator_0/un6lto15_1 )
        , .B(\modulator_0/un6lt15 ), .C(
        \modulator_0/output_signal_1_sqmuxa_0 ), .Y(
        \modulator_0/output_signal_1_sqmuxa_0_0 ));
    DFN1E1P0 \data_source_0/tag_data_buf_5[2]  (.D(
        \data_source_0/tag_data_buf_5_4[2] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_5[2]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_8[8]  (.A(
        \data_source_0/N_729 ), .B(\data_source_0/N_1189 ), .C(
        \data_source_0/N_949 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[8] ));
    OR3 \data_source_0/tag_control_sig_RNO_3[13]  (.A(
        \data_source_0/N_1223 ), .B(\data_source_0/N_1224 ), .C(
        \data_source_0/N_1028 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[13] ));
    MX2 \switching_circuit_0/out_signal_switch_1[3]  (.A(
        \switching_circuit_0/un30_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un33_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[3] ));
    DFN1E1C0 \data_source_0/tag_data_buf_19[2]  (.D(
        \data_source_0/tag_data_buf_19_4[2] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_19[2]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_8[13]  (.A(
        \data_source_0/N_996_1 ), .B(\data_source_0/N_1204 ), .C(
        \data_source_0/N_1024 ), .Y(
        \data_source_0/tag_control_sig_2_0_9[13] ));
    NOR2B \data_source_0/tag_data_buf_6_RNO[4]  (.A(
        \data_source_0/tag_data_buf_6[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_6_4[4] ));
    DFN1E1C0 \data_source_0/tag_data_buf_19[3]  (.D(
        \data_source_0/tag_data_buf_19_4[3] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_19[3]_net_1 ));
    IOIN_IB \trigger_signal_pad/U0/U1  (.YIN(
        \trigger_signal_pad/U0/NET1 ), .Y(trigger_signal_c));
    OA1 \data_source_0/data_index_RNIR3731[6]  (.A(
        \data_source_0/N_1155 ), .B(\data_source_0/N_1171 ), .C(
        \data_source_0/N_1134 ), .Y(\data_source_0/N_1245 ));
    AO1 \data_source_0/tag_control_sig_RNO_19[5]  (.A(
        \data_source_0/N_804 ), .B(\data_source_0/N_1191 ), .C(
        \data_source_0/N_902 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[5] ));
    DFN1E1C0 \data_source_0/output_data[19]  (.D(
        \data_source_0/output_data_23[19] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[19] ));
    OR3 \data_source_0/tag_control_sig_RNO_1[14]  (.A(
        \data_source_0/N_1044 ), .B(\data_source_0/N_1041 ), .C(
        \data_source_0/tag_control_sig_2_0_6[14] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[14] ));
    NOR2B \data_source_0/data_index_RNI9K6D_0[6]  (.A(
        \data_source_0/N_1133 ), .B(
        \data_source_0/data_index[6]_net_1 ), .Y(
        \data_source_0/N_1154 ));
    NOR2B \data_source_0/tag_data_buf_20_RNO[7]  (.A(
        \data_source_0/tag_data_buf_20[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_20_4[7] ));
    NOR2B \data_source_0/tag_data_buf_1_RNO[1]  (.A(
        \data_source_0/tag_data_buf_1[0]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_1_4[1] ));
    OR3 \data_source_0/tag_control_sig_RNO[0]  (.A(
        \data_source_0/tag_control_sig_2_0_13[0] ), .B(
        \data_source_0/tag_control_sig_2_0_12[0] ), .C(
        \data_source_0/tag_control_sig_2_0_14[0] ), .Y(
        \data_source_0/tag_control_sig_2[0] ));
    NOR2B \data_source_0/tag_control_sig_RNO_7[2]  (.A(
        \data_source_0/N_1192 ), .B(\data_source_0/N_1161 ), .Y(
        \data_source_0/N_862 ));
    OR3 \data_source_0/tag_control_sig_RNO[11]  (.A(
        \data_source_0/tag_control_sig_2_0_16[11] ), .B(
        \data_source_0/tag_control_sig_2_0_15[11] ), .C(
        \data_source_0/tag_control_sig_2_0_17[11] ), .Y(
        \data_source_0/tag_control_sig_2[11] ));
    NOR2B \data_source_0/tag_data_buf_8_RNI0GBJ[7]  (.A(
        \data_source_0/tag_data_buf_8[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[7] ));
    NOR3B \data_source_0/data_index_0_RNI1NTK[7]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/N_1141 ), .C(
        \data_source_0/data_index_0[7]_net_1 ), .Y(
        \data_source_0/N_1198 ));
    AO1 \data_source_0/tag_control_sig_RNO_4[19]  (.A(
        \data_source_0/N_1187 ), .B(\data_source_0/N_1161 ), .C(
        \data_source_0/N_860 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[19] ));
    NOR2A \data_source_0/data_index_RNIASP8[4]  (.A(
        \data_source_0/data_index[4]_net_1 ), .B(
        \data_source_0/data_index[6]_net_1 ), .Y(
        \data_source_0/N_1208 ));
    NOR3C \data_source_0/tag_control_sig_RNO_6[18]  (.A(
        \data_source_0/tag_control_sig_1_3[649] ), .B(
        \data_source_0/N_1148 ), .C(\data_source_0/N_1182 ), .Y(
        \data_source_0/N_1110 ));
    DFN1E1P0 \data_source_0/tag_data_buf_2[1]  (.D(
        \data_source_0/tag_data_buf_2_4[1] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_2[1]_net_1 ));
    NOR2A \data_source_0/data_index_RNI9K6D[3]  (.A(
        \data_source_0/N_703_i ), .B(
        \data_source_0/data_index[3]_net_1 ), .Y(
        \data_source_0/N_1234 ));
    NOR2B \data_source_0/tag_data_buf_15_RNO[5]  (.A(
        \data_source_0/tag_data_buf_15[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_15_4[5] ));
    OR3 \data_source_0/tag_control_sig_RNO_2[14]  (.A(
        \data_source_0/tag_control_sig_2_0_5[14] ), .B(
        \data_source_0/tag_control_sig_2_0_4[14] ), .C(
        \data_source_0/tag_control_sig_2_0_10[14] ), .Y(
        \data_source_0/tag_control_sig_2_0_14[14] ));
    XOR2 \main_clock_0/un5_counter_1_I_14  (.A(\main_clock_0/N_4 ), .B(
        \main_clock_0/counter[5]_net_1 ), .Y(\main_clock_0/I_14_0 ));
    NOR3C \data_source_0/tag_control_sig_RNO_17[10]  (.A(
        \data_source_0/data_index[3]_net_1 ), .B(
        \data_source_0/N_1145 ), .C(
        \data_source_0/tag_control_sig_2_0_a20_4_0[10] ), .Y(
        \data_source_0/N_978 ));
    NOR2B \data_source_0/tag_control_sig_RNO_15[5]  (.A(
        \data_source_0/N_1137 ), .B(\data_source_0/N_1174 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_3_0[5] ));
    AO1A \data_source_0/tag_control_sig_RNO_19[16]  (.A(
        \data_source_0/N_759 ), .B(
        \data_source_0/tag_control_sig_2_0_a20_4_0[16] ), .C(
        \data_source_0/N_1082 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[16] ));
    AO1 \data_source_0/tag_control_sig_RNO_10[11]  (.A(
        \data_source_0/N_1202 ), .B(\data_source_0/N_1161 ), .C(
        \data_source_0/N_1000 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[11] ));
    DFN1E1C0 \data_source_0/output_data[16]  (.D(
        \data_source_0/output_data_23[16] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[16] ));
    AO1 \data_source_0/tag_control_sig_RNO_18[0]  (.A(
        \data_source_0/N_1190 ), .B(\data_source_0/N_1184 ), .C(
        \data_source_0/N_818 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[0] ));
    IOTRI_OB_EB \output_signal_pad[3]/U0/U1  (.D(\output_signal_c[3] ), 
        .E(VCC), .DOUT(\output_signal_pad[3]/U0/NET1 ), .EOUT(
        \output_signal_pad[3]/U0/NET2 ));
    XA1 \modulator_0/clock_counter_RNO[13]  (.A(
        \modulator_0/clock_counter_c12 ), .B(
        \modulator_0/clock_counter[13]_net_1 ), .C(AND2_0_Y), .Y(
        \modulator_0/clock_counter_n13 ));
    NOR2B \data_source_0/tag_data_buf_13_RNO[6]  (.A(
        \data_source_0/tag_data_buf_13[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_13_4[6] ));
    NOR2B \data_source_0/data_index_RNIRO0M_2[7]  (.A(
        \data_source_0/N_1138 ), .B(\data_source_0/N_1143 ), .Y(
        \data_source_0/N_1176 ));
    XA1A \switching_circuit_0/un73_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[7] ), 
        .C(\data_source_0_tag_control_sig[7] ), .Y(
        \switching_circuit_0/un73_out_signal_switch_0_net_1 ));
    AOI1D \data_source_0/tag_control_sig_RNO_4[12]  (.A(
        \data_source_0/N_1200 ), .B(\data_source_0/N_1199 ), .C(
        \data_source_0/N_1180 ), .Y(
        \data_source_0/tag_control_sig_RNO_4[12]_net_1 ));
    DFN1C0 \main_clock_0/counter[3]  (.D(\main_clock_0/I_9_0 ), .CLK(
        GLA), .CLR(reset_c), .Q(\main_clock_0/counter[3]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_7[6]  (.D(
        \data_source_0/tag_data_buf_7_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_7[6]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_2[7]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_6_0[7] ), .B(
        \data_source_0/N_1191 ), .C(\data_source_0/N_935 ), .Y(
        \data_source_0/tag_control_sig_2_0_6[7] ));
    OR3 \modulator_0/output_signal_RNO_10  (.A(\modulator_0/un6lto9 ), 
        .B(\modulator_0/clock_counter[15]_net_1 ), .C(
        \modulator_0/un6lto10 ), .Y(\modulator_0/un5lto15_3 ));
    DFN1E1P0 \data_source_0/tag_data_buf_11[3]  (.D(
        \data_source_0/tag_data_buf_11_4[3] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_11[3]_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_16[8]  (.A(
        \data_source_0/data_index_0[7]_net_1 ), .B(
        \data_source_0/N_1135 ), .C(
        \data_source_0/tag_control_sig_2_0_a20_6_0[8] ), .Y(
        \data_source_0/N_949 ));
    NOR2B \data_source_0/data_index_0_RNIJ6UA1_1[7]  (.A(
        \data_source_0/N_1191 ), .B(\data_source_0/N_1185 ), .Y(
        \data_source_0/N_832 ));
    NOR3A \data_source_0/tag_control_sig_RNO_12[5]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/data_index_0[7]_net_1 ), .C(
        \data_source_0/data_index[3]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_1_1[5] ));
    XA1 \modulator_0/counter_RNO[5]  (.A(
        \modulator_0/counter[5]_net_1 ), .B(\modulator_0/counter_45_0 )
        , .C(\modulator_0/counter_0_sqmuxa ), .Y(
        \modulator_0/counter_n5 ));
    DFN1E1C0 \data_source_0/tag_data_buf_5[7]  (.D(
        \data_source_0/tag_data_buf_5_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_5[7]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_8[9]  (.A(
        \data_source_0/N_1192 ), .B(\data_source_0/N_1182 ), .C(
        \data_source_0/N_961 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[9] ));
    DFN1E1 \data_source_0/tag_control_sig[2]  (.D(
        \data_source_0/tag_control_sig_2[2] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[2] ));
    NOR2B \data_source_0/tag_data_buf_1_RNO[4]  (.A(
        \data_source_0/tag_data_buf_1[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_1_4[4] ));
    NOR2B \data_source_0/data_index_RNIO37D[7]  (.A(
        \data_source_0/N_1139 ), .B(
        \data_source_0/data_index[7]_net_1 ), .Y(
        \data_source_0/N_1237 ));
    OR2 \data_source_0/counter_RNI2OR61[3]  (.A(
        \data_source_0/counter_i_0[3] ), .B(\data_source_0/N_32 ), .Y(
        \data_source_0/N_33 ));
    XA1A \data_source_0/counter_RNO[10]  (.A(\data_source_0/N_39 ), .B(
        \data_source_0/counter[10]_net_1 ), .C(
        modulator_0_output_signal), .Y(\data_source_0/counter_n10 ));
    MX2 \switching_circuit_0/out_signal_switch_1[6]  (.A(
        \switching_circuit_0/un60_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un63_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[6] ));
    NOR2B \data_source_0/tag_data_buf_2_RNO[2]  (.A(
        \data_source_0/tag_data_buf_2[1]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_2_4[2] ));
    NOR2A \data_source_0/data_index_RNI7PP8_1[1]  (.A(
        \data_source_0/data_index[6]_net_1 ), .B(
        \data_source_0/data_index[1]_net_1 ), .Y(
        \data_source_0/N_1137 ));
    DFN1E1P0 \data_source_0/tag_data_buf_4[2]  (.D(
        \data_source_0/tag_data_buf_4_4[2] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_4[2]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_9[2]  (.A(
        \data_source_0/N_729 ), .B(\data_source_0/N_1209 ), .C(
        \data_source_0/N_849 ), .Y(
        \data_source_0/tag_control_sig_2_0_2[2] ));
    OR3 \data_source_0/tag_control_sig_RNO_1[6]  (.A(
        \data_source_0/N_915 ), .B(\data_source_0/N_914 ), .C(
        \data_source_0/tag_control_sig_2_0_3[6] ), .Y(
        \data_source_0/tag_control_sig_2_0_10[6] ));
    XA1 \modulator_0/clock_counter_RNO[4]  (.A(
        \modulator_0/clock_counter[4]_net_1 ), .B(
        \modulator_0/clock_counter_c3 ), .C(AND2_0_Y), .Y(
        \modulator_0/clock_counter_n4 ));
    NOR2B \data_source_0/tag_control_sig_RNO_6[2]  (.A(
        \data_source_0/N_1197 ), .B(\data_source_0/N_1163 ), .Y(
        \data_source_0/N_863 ));
    NOR2B \data_source_0/data_index_RNI46K71_0[5]  (.A(
        \data_source_0/N_1191 ), .B(\data_source_0/N_1162 ), .Y(
        \data_source_0/N_1028 ));
    DFN1E1C0 \data_source_0/tag_data_buf_12[7]  (.D(
        \data_source_0/tag_data_buf_12_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_12[7]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_11[16]  (.A(
        \data_source_0/tag_control_sig_RNO_17[16]_net_1 ), .B(
        \data_source_0/N_1073 ), .C(
        \data_source_0/tag_control_sig_2_0_7[16] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[16] ));
    OR2 \data_source_0/tag_control_sig_RNO_23[5]  (.A(
        \data_source_0/N_1173 ), .B(\data_source_0/N_1174 ), .Y(
        \data_source_0/N_804 ));
    NOR2B \data_source_0/tag_control_sig_RNO_11[6]  (.A(
        \data_source_0/N_1140 ), .B(\data_source_0/N_1176 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_3_0[6] ));
    DFN1E1C0 \data_source_0/tag_data_buf_14[6]  (.D(
        \data_source_0/tag_data_buf_14_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_14[6]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_2_RNO[3]  (.A(
        \data_source_0/tag_data_buf_2[2]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_2_4[3] ));
    NOR2B \data_source_0/tag_control_sig_RNO_20[18]  (.A(
        \data_source_0/N_1192 ), .B(\data_source_0/N_1160 ), .Y(
        \data_source_0/N_1109 ));
    NOR2B \data_source_0/tag_control_sig_RNO_19[17]  (.A(
        \data_source_0/N_1187 ), .B(\data_source_0/N_1178 ), .Y(
        \data_source_0/N_1098 ));
    IOTRI_OB_EB \output_signal_pad[16]/U0/U1  (.D(
        \output_signal_c[16] ), .E(VCC), .DOUT(
        \output_signal_pad[16]/U0/NET1 ), .EOUT(
        \output_signal_pad[16]/U0/NET2 ));
    NOR2B \data_source_0/tag_control_sig_RNO_19[3]  (.A(
        \data_source_0/N_1205 ), .B(\data_source_0/N_1142 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_9_0[3] ));
    OR3 \data_source_0/tag_control_sig_RNO_0[19]  (.A(
        \data_source_0/tag_control_sig_RNO_3[19]_net_1 ), .B(
        \data_source_0/N_1010 ), .C(
        \data_source_0/tag_control_sig_2_0_7[19] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[19] ));
    XA1A \switching_circuit_0/un193_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[19] ), 
        .C(\data_source_0_tag_control_sig[19] ), .Y(
        \switching_circuit_0/un193_out_signal_switch_0_net_1 ));
    IOIN_IB \clock_pad/U0/U1  (.YIN(\clock_pad/U0/NET1 ), .Y(clock_c));
    NOR2A \data_source_0/data_index_RNIJNJH[7]  (.A(
        \data_source_0/N_1159 ), .B(
        \data_source_0/data_index[7]_net_1 ), .Y(
        \data_source_0/N_996_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_5[4]  (.D(
        \data_source_0/tag_data_buf_5_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_5[4]_net_1 ));
    NOR2B \data_source_0/data_index_RNI9K6D[2]  (.A(
        \data_source_0/N_1137 ), .B(
        \data_source_0/data_index[2]_net_1 ), .Y(
        \data_source_0/N_1157 ));
    NOR2B \data_source_0/tag_control_sig_RNO_16[5]  (.A(
        \data_source_0/N_1210 ), .B(\data_source_0/N_1162 ), .Y(
        \data_source_0/N_911 ));
    AO1A \data_source_0/tag_control_sig_RNO_17[1]  (.A(
        \data_source_0/N_759 ), .B(
        \data_source_0/tag_control_sig_2_0_a20_6_0[1] ), .C(
        \data_source_0/N_835 ), .Y(
        \data_source_0/tag_control_sig_2_0_2[1] ));
    DFN1E1P0 \data_source_0/tag_data_buf_10[3]  (.D(
        \data_source_0/tag_data_buf_10_4[3] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_10[3]_net_1 ));
    NOR3C \data_source_0/tag_control_sig_RNO_4[16]  (.A(
        \data_source_0/N_1140 ), .B(\data_source_0/N_1154 ), .C(
        \data_source_0/N_1184 ), .Y(\data_source_0/N_1083 ));
    OR3 \data_source_0/tag_control_sig_RNO_0[12]  (.A(
        \data_source_0/N_1015 ), .B(
        \data_source_0/tag_control_sig_RNO_4[12]_net_1 ), .C(
        \data_source_0/tag_control_sig_2_0_7[12] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[12] ));
    AX1C \main_clock_0/un5_counter_1_I_7  (.A(
        \main_clock_0/counter[1]_net_1 ), .B(
        \main_clock_0/counter[0]_net_1 ), .C(
        \main_clock_0/counter[2]_net_1 ), .Y(\main_clock_0/I_7_0 ));
    NOR2B \data_source_0/tag_control_sig_RNO_12[8]  (.A(
        \data_source_0/N_1206 ), .B(\data_source_0/N_1177 ), .Y(
        \data_source_0/N_954 ));
    NOR3C \data_source_0/data_index_RNI4D731[0]  (.A(
        \data_source_0/tag_control_sig_1_649_1 ), .B(
        \data_source_0/tag_control_sig_1_649_0 ), .C(
        \data_source_0/tag_control_sig_1_649_5 ), .Y(
        \data_source_0/tag_control_sig_1_649_6 ));
    OR3 \data_source_0/tag_control_sig_RNO_1[3]  (.A(
        \data_source_0/N_873 ), .B(\data_source_0/N_872 ), .C(
        \data_source_0/tag_control_sig_2_0_1[3] ), .Y(
        \data_source_0/tag_control_sig_2_0_9[3] ));
    AO1 \data_source_0/tag_control_sig_RNO_4[11]  (.A(
        \data_source_0/N_1189 ), .B(\data_source_0/N_1185 ), .C(
        \data_source_0/N_995 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[11] ));
    OA1 \data_source_0/tag_control_sig_RNO_13[2]  (.A(
        \data_source_0/N_1244 ), .B(\data_source_0/N_1235 ), .C(
        \data_source_0/N_1193 ), .Y(
        \data_source_0/tag_control_sig_RNO_13[2]_net_1 ));
    NOR2 \data_source_0/data_index_RNIG2Q8[9]  (.A(
        \data_source_0/data_index[9]_net_1 ), .B(
        \data_source_0/data_index[7]_net_1 ), .Y(
        \data_source_0/N_1240 ));
    NOR2B \data_source_0/tag_control_sig_RNO_6[5]  (.A(
        \data_source_0/N_1226 ), .B(\data_source_0/N_1159 ), .Y(
        \data_source_0/N_907 ));
    AOI1D \data_source_0/tag_control_sig_RNO_5[4]  (.A(
        \data_source_0/N_1184 ), .B(\data_source_0/N_1175 ), .C(
        \data_source_0/N_1190 ), .Y(\data_source_0/N_881 ));
    NOR2A \modulator_0/counter_RNIBT613[4]  (.A(AND2_0_Y), .B(
        \modulator_0/counter19 ), .Y(\modulator_0/counter_0_sqmuxa ));
    NOR2B \data_source_0/tag_data_buf_4_RNO[7]  (.A(
        \data_source_0/tag_data_buf_4[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_4_4[7] ));
    DFN1E1C0 \data_source_0/tag_data_buf_12[1]  (.D(
        \data_source_0/tag_data_buf_12_4[1] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_12[1]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_3_RNO[5]  (.A(
        \data_source_0/tag_data_buf_3[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_3_4[5] ));
    OR3 \data_source_0/tag_control_sig_RNO_11[17]  (.A(
        \data_source_0/N_1096 ), .B(\data_source_0/N_1094 ), .C(
        \data_source_0/tag_control_sig_2_0_5[17] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[17] ));
    NOR3A \data_source_0/tag_control_sig_RNO_6[8]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_10_0[8] ), .B(
        \data_source_0/data_index_0[7]_net_1 ), .C(
        \data_source_0/data_index[8]_net_1 ), .Y(\data_source_0/N_953 )
        );
    OR3 \data_source_0/tag_control_sig_RNO[15]  (.A(
        \data_source_0/tag_control_sig_2_0_14[15] ), .B(
        \data_source_0/tag_control_sig_2_0_13[15] ), .C(
        \data_source_0/tag_control_sig_2_0_15[15] ), .Y(
        \data_source_0/tag_control_sig_2[15] ));
    DFN1E1C0 \modulator_0/clock_counter[6]  (.D(
        \modulator_0/clock_counter_n6 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/un5lto6 ));
    OR2A \data_source_0/counter_RNI4GC23[11]  (.A(
        \data_source_0/counter[11]_net_1 ), .B(\data_source_0/N_40 ), 
        .Y(\data_source_0/N_41 ));
    AND3 \data_source_0/un3_data_index_I_8  (.A(
        \data_source_0/data_index[0]_net_1 ), .B(
        \data_source_0/data_index[1]_net_1 ), .C(
        \data_source_0/data_index[2]_net_1 ), .Y(\data_source_0/N_8 ));
    NOR2B \data_source_0/tag_data_buf_19_RNO[3]  (.A(
        \data_source_0/tag_data_buf_19[2]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_19_4[3] ));
    XA1A \data_source_0/counter_RNO[15]  (.A(\data_source_0/N_44 ), .B(
        \data_source_0/counter[15]_net_1 ), .C(
        modulator_0_output_signal), .Y(\data_source_0/counter_n15 ));
    DFN1P0 \data_source_0/counter[6]  (.D(\data_source_0/N_16 ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .Q(
        \data_source_0/counter_i_0[6] ));
    DFN1E1C0 \data_source_0/tag_data_buf_17[1]  (.D(
        \data_source_0/tag_data_buf_17_4[1] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_17[1]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_15[14]  (.A(
        \data_source_0/N_1173 ), .B(\data_source_0/N_1198 ), .C(
        \data_source_0/N_1186 ), .Y(\data_source_0/N_802 ));
    NOR2B \data_source_0/tag_control_sig_RNO_7[0]  (.A(
        \data_source_0/N_1199 ), .B(\data_source_0/N_1161 ), .Y(
        \data_source_0/N_825 ));
    AOI1B \data_source_0/data_index_RNIODII2[4]  (.A(
        \data_source_0/tag_control_sig_1_649_6 ), .B(
        \data_source_0/tag_control_sig_1_3[649] ), .C(
        \data_source_0/I_20 ), .Y(\data_source_0/data_index_3[7] ));
    DFN1E1C0 \data_source_0/tag_data_buf_20[5]  (.D(
        \data_source_0/tag_data_buf_20_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_20[5]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_3[15]  (.A(
        \data_source_0/N_778 ), .B(\data_source_0/N_1173 ), .C(
        \data_source_0/N_1058 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[15] ));
    NOR2A \data_source_0/tag_control_sig_1_sqmuxa  (.A(reset_c), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_10[12]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_1_1[12] ), .B(
        \data_source_0/tag_control_sig_2_0_a20_1_0[12] ), .C(
        \data_source_0/N_835 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[12] ));
    NOR2B \data_source_0/tag_data_buf_7_RNO[3]  (.A(
        \data_source_0/tag_data_buf_7[2]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_7_4[3] ));
    AO1 \data_source_0/tag_control_sig_RNO_8[15]  (.A(
        \data_source_0/N_1225 ), .B(\data_source_0/N_1177 ), .C(
        \data_source_0/N_1063 ), .Y(
        \data_source_0/tag_control_sig_2_0_8[15] ));
    NOR2B \data_source_0/data_index_RNIIF0M_8[6]  (.A(
        \data_source_0/N_1156 ), .B(\data_source_0/N_1154 ), .Y(
        \data_source_0/N_1226 ));
    XA1 \modulator_0/clock_counter_RNO[6]  (.A(
        \modulator_0/clock_counter_c5 ), .B(\modulator_0/un5lto6 ), .C(
        AND2_0_Y), .Y(\modulator_0/clock_counter_n6 ));
    DFN1E1C0 \data_source_0/tag_data_buf_13[5]  (.D(
        \data_source_0/tag_data_buf_13_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_13[5]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_1[9]  (.A(
        \data_source_0/N_962 ), .B(\data_source_0/N_969 ), .C(
        \data_source_0/tag_control_sig_2_0_7[9] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[9] ));
    NOR2B \data_source_0/tag_data_buf_3_RNO[7]  (.A(
        \data_source_0/tag_data_buf_3[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_3_4[7] ));
    DFN1E1 \data_source_0/tag_control_sig[6]  (.D(
        \data_source_0/tag_control_sig_2[6] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[6] ));
    NOR3B \data_source_0/data_index_0_RNI1NTK_0[7]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/N_1138 ), .C(
        \data_source_0/data_index_0[7]_net_1 ), .Y(
        \data_source_0/N_1180 ));
    IOTRI_OB_EB \output_signal_pad[19]/U0/U1  (.D(
        \output_signal_c[19] ), .E(VCC), .DOUT(
        \output_signal_pad[19]/U0/NET1 ), .EOUT(
        \output_signal_pad[19]/U0/NET2 ));
    AO1 \data_source_0/tag_control_sig_RNO_5[19]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_1_0[19] ), .B(
        \data_source_0/N_868_1 ), .C(\data_source_0/N_1120 ), .Y(
        \data_source_0/tag_control_sig_2_0_4[19] ));
    NOR2B \data_source_0/tag_control_sig_RNO_22[5]  (.A(
        \data_source_0/N_1138 ), .B(
        \data_source_0/data_index[8]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_10_0[5] ));
    NOR2B \data_source_0/data_index_RNIBM6D[1]  (.A(
        \data_source_0/N_1208 ), .B(
        \data_source_0/data_index[1]_net_1 ), .Y(
        \data_source_0/N_1232 ));
    OR3 \data_source_0/tag_control_sig_RNO_9[12]  (.A(
        \data_source_0/N_921 ), .B(\data_source_0/N_1218 ), .C(
        \data_source_0/N_1007 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[12] ));
    DFN1E1C0 \modulator_0/output_signal  (.D(
        \modulator_0/output_signal_1_sqmuxa_0_0 ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \modulator_0/clock_countere ), .Q(
        \modulator_0/output_signal_i ));
    OR3 \data_source_0/tag_control_sig_RNO_0[16]  (.A(
        \data_source_0/N_1080 ), .B(\data_source_0/N_1083 ), .C(
        \data_source_0/tag_control_sig_2_0_2[16] ), .Y(
        \data_source_0/tag_control_sig_2_0_9[16] ));
    OR2A \data_source_0/counter_RNI9Q9Q1[5]  (.A(
        \data_source_0/counter[5]_net_1 ), .B(\data_source_0/N_34 ), 
        .Y(\data_source_0/N_35 ));
    DFN1C0 \main_clock_0/counter[5]  (.D(\main_clock_0/I_14_0 ), .CLK(
        GLA), .CLR(reset_c), .Q(\main_clock_0/counter[5]_net_1 ));
    NOR2B \switching_circuit_0/un20_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[2] ), .B(main_clock_0_clock_out)
        , .Y(\switching_circuit_0/un20_out_signal_switch_0_net_1 ));
    NOR3B \data_source_0/tag_control_sig_RNO_20[12]  (.A(
        \data_source_0/N_1157 ), .B(\data_source_0/N_1163 ), .C(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/N_1013 ));
    NOR2B \data_source_0/tag_data_buf_1_RNO[5]  (.A(
        \data_source_0/tag_data_buf_1[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_1_4[5] ));
    OR2A \data_source_0/tag_data_buf_11_RNO[3]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_11[2]_net_1 ), .Y(
        \data_source_0/tag_data_buf_11_4[3] ));
    NOR3C \data_source_0/tag_control_sig_RNO_20[15]  (.A(
        \data_source_0/N_1133 ), .B(\data_source_0/N_1151 ), .C(
        \data_source_0/N_1179 ), .Y(\data_source_0/N_1066 ));
    OR3 \data_source_0/tag_control_sig_RNO_0[11]  (.A(
        \data_source_0/tag_control_sig_2_0_2[11] ), .B(
        \data_source_0/tag_control_sig_2_0_1[11] ), .C(
        \data_source_0/tag_control_sig_2_0_12[11] ), .Y(
        \data_source_0/tag_control_sig_2_0_16[11] ));
    DFN1E1P0 \data_source_0/tag_data_buf_8[3]  (.D(
        \data_source_0/tag_data_buf_8_4[3] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_8[3]_net_1 ));
    OR2A \data_source_0/tag_data_buf_18_RNO[1]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_18[0]_net_1 ), .Y(
        \data_source_0/tag_data_buf_18_4[1] ));
    OR3 \data_source_0/tag_control_sig_RNO_1[5]  (.A(
        \data_source_0/N_907 ), .B(\data_source_0/N_909 ), .C(
        \data_source_0/tag_control_sig_2_0_6[5] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[5] ));
    AO1 \data_source_0/tag_control_sig_RNO_10[9]  (.A(
        \data_source_0/N_777 ), .B(\data_source_0/N_1159 ), .C(
        \data_source_0/N_957 ), .Y(
        \data_source_0/tag_control_sig_2_0_2[9] ));
    AND3 \main_clock_0/un5_counter_1_I_13  (.A(
        \main_clock_0/DWACT_FINC_E[0] ), .B(
        \main_clock_0/counter[3]_net_1 ), .C(
        \main_clock_0/counter[4]_net_1 ), .Y(\main_clock_0/N_4 ));
    AX1C \main_clock_0/un5_counter_1_I_12  (.A(
        \main_clock_0/counter[3]_net_1 ), .B(
        \main_clock_0/DWACT_FINC_E[0] ), .C(
        \main_clock_0/counter[4]_net_1 ), .Y(\main_clock_0/I_12_0 ));
    AO1 \data_source_0/tag_control_sig_RNO_5[12]  (.A(
        \data_source_0/N_1209 ), .B(\data_source_0/N_1160 ), .C(
        \data_source_0/N_1014 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[12] ));
    NOR2B \data_source_0/data_index_RNIIF0M_0[2]  (.A(
        \data_source_0/N_1157 ), .B(\data_source_0/N_1140 ), .Y(
        \data_source_0/N_1202 ));
    NOR2B \modulator_0/clock_counter_RNID686[4]  (.A(
        \modulator_0/clock_counter_c3 ), .B(
        \modulator_0/clock_counter[4]_net_1 ), .Y(
        \modulator_0/clock_counter_c4 ));
    CLKINT \modulator_0/output_signal_RNI2QGD  (.A(
        \modulator_0/output_signal_i ), .Y(modulator_0_output_signal));
    NOR2B \data_source_0/data_index_RNICN6D[9]  (.A(
        \data_source_0/data_index[9]_net_1 ), .B(
        \data_source_0/N_1132 ), .Y(\data_source_0/N_1159 ));
    XA1 \modulator_0/clock_counter_RNO[9]  (.A(
        \modulator_0/clock_counter_c8 ), .B(\modulator_0/un6lto9 ), .C(
        AND2_0_Y), .Y(\modulator_0/clock_counter_n9 ));
    CLKINT \data_source_0/counter_RNIK0AI3_0[1]  (.A(
        \data_source_0/counter_RNIK0AI3[1]_net_1 ), .Y(
        \data_source_0/N_29 ));
    DFN1C0 \main_clock_0/counter[2]  (.D(\main_clock_0/I_7_0 ), .CLK(
        GLA), .CLR(reset_c), .Q(\main_clock_0/counter[2]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_18_RNIHCFR[7]  (.A(
        \data_source_0/tag_data_buf_18[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[17] ));
    NOR2B \data_source_0/data_index_RNIF1Q8[7]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/data_index[7]_net_1 ), .Y(
        \data_source_0/N_1144 ));
    NOR2A \data_source_0/data_index_RNIFQ6D[6]  (.A(
        \data_source_0/N_1140 ), .B(
        \data_source_0/data_index[6]_net_1 ), .Y(
        \data_source_0/N_1158 ));
    NOR2A \data_source_0/data_index_RNI9K6D_0[2]  (.A(
        \data_source_0/N_1137 ), .B(
        \data_source_0/data_index[2]_net_1 ), .Y(
        \data_source_0/N_1155 ));
    NOR3A \modulator_0/counter_RNIUHHV1[5]  (.A(
        \modulator_0/counter19_3 ), .B(\modulator_0/counter[4]_net_1 ), 
        .C(\modulator_0/counter[5]_net_1 ), .Y(
        \modulator_0/counter23_2 ));
    NOR2B \data_source_0/tag_control_sig_RNO_17[14]  (.A(
        \data_source_0/N_1225 ), .B(\data_source_0/N_1198 ), .Y(
        \data_source_0/N_1050 ));
    DFN1E1P0 \data_source_0/tag_data_buf_18[1]  (.D(
        \data_source_0/tag_data_buf_18_4[1] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_18[1]_net_1 ));
    DFN1E1P0 \data_source_0/tag_data_buf_3[1]  (.D(
        \data_source_0/tag_data_buf_3_4[1] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_3[1]_net_1 ));
    NOR2B \data_source_0/data_index_RNI9RP8[4]  (.A(
        \data_source_0/data_index[4]_net_1 ), .B(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/N_1134 ));
    NOR2A \data_source_0/data_index_RNI9RP8_1[4]  (.A(
        \data_source_0/data_index[4]_net_1 ), .B(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/N_1140 ));
    NOR2B \data_source_0/tag_control_sig_RNO_22[19]  (.A(
        \data_source_0/N_1197 ), .B(\data_source_0/N_1160 ), .Y(
        \data_source_0/N_1122 ));
    NOR2B \data_source_0/tag_control_sig_RNO_24[17]  (.A(
        \data_source_0/N_1183 ), .B(\data_source_0/N_1163 ), .Y(
        \data_source_0/N_1101 ));
    OR2 \data_source_0/data_index_RNI4V0C1[6]  (.A(
        \data_source_0/N_1188 ), .B(\data_source_0/N_1190 ), .Y(
        \data_source_0/N_766 ));
    OR2 \modulator_0/output_signal_RNO_8  (.A(
        \modulator_0/clock_counter[14]_net_1 ), .B(
        \modulator_0/clock_counter[13]_net_1 ), .Y(
        \modulator_0/un5lto15_2 ));
    OR3 \data_source_0/tag_control_sig_RNO_0[0]  (.A(
        \data_source_0/tag_control_sig_2_0_1[0] ), .B(
        \data_source_0/tag_control_sig_2_0_0[0] ), .C(
        \data_source_0/tag_control_sig_2_0_8[0] ), .Y(
        \data_source_0/tag_control_sig_2_0_13[0] ));
    OR2A \data_source_0/tag_data_buf_15_RNO[1]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_15[0]_net_1 ), .Y(
        \data_source_0/tag_data_buf_15_4[1] ));
    DFN1E1C0 \data_source_0/tag_data_buf_10[0]  (.D(
        \data_source_0/output_data_23[9] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_10[0]_net_1 ));
    NOR3B \data_source_0/tag_control_sig_RNO_22[16]  (.A(
        \data_source_0/N_1237 ), .B(
        \data_source_0/tag_control_sig_2_0_a20_9_2[16] ), .C(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/N_1082 ));
    DFN1E1C0 \data_source_0/tag_data_buf_16[5]  (.D(
        \data_source_0/tag_data_buf_16_4[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_16[5]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_22[8]  (.A(
        \data_source_0/N_1208 ), .B(\data_source_0/N_1173 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_4_0[8] ));
    NOR3C \data_source_0/tag_control_sig_RNO_15[18]  (.A(
        \data_source_0/N_1133 ), .B(\data_source_0/N_1151 ), .C(
        \data_source_0/N_1184 ), .Y(\data_source_0/N_1115 ));
    XAI1 \data_source_0/counter_RNO[4]  (.A(\data_source_0/N_33 ), .B(
        \data_source_0/counter_i_0[4] ), .C(modulator_0_output_signal), 
        .Y(\data_source_0/N_20 ));
    NOR3B \data_source_0/tag_control_sig_RNO_23[16]  (.A(
        \data_source_0/N_1149 ), .B(\data_source_0/N_1141 ), .C(
        \data_source_0/data_index[6]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_9_2[16] ));
    DFN1E1 \data_source_0/tag_control_sig[3]  (.D(
        \data_source_0/tag_control_sig_2[3] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[3] ));
    NOR2B \data_source_0/tag_control_sig_RNO_10[4]  (.A(
        \data_source_0/N_1136 ), .B(\data_source_0/N_1134 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_8_0[4] ));
    NOR2B \data_source_0/data_index_RNIIF0M_4[6]  (.A(
        \data_source_0/N_1158 ), .B(\data_source_0/N_1133 ), .Y(
        \data_source_0/N_1192 ));
    NOR2A \data_source_0/data_index_RNIH3Q8[9]  (.A(
        \data_source_0/data_index[9]_net_1 ), .B(
        \data_source_0/data_index[8]_net_1 ), .Y(
        \data_source_0/tag_control_sig_1_649_0 ));
    DFN1E1C0 \data_source_0/tag_data_buf_14[7]  (.D(
        \data_source_0/tag_data_buf_14_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_14[7]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_9[16]  (.A(
        \data_source_0/N_1202 ), .B(\data_source_0/N_1175 ), .C(
        \data_source_0/N_1078 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[16] ));
    NOR2B \data_source_0/tag_control_sig_RNO_18[19]  (.A(
        \data_source_0/N_701_i ), .B(\data_source_0/N_1174 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_2_0[19] ));
    DFN1E1P0 \data_source_0/tag_data_buf_13[3]  (.D(
        \data_source_0/tag_data_buf_13_4[3] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_13[3]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_9[11]  (.A(
        \data_source_0/N_996_1 ), .B(\data_source_0/N_1187 ), .C(
        \data_source_0/N_904 ), .Y(
        \data_source_0/tag_control_sig_2_0_6[11] ));
    OA1 \data_source_0/tag_control_sig_RNO_8[5]  (.A(
        \data_source_0/N_1189 ), .B(\data_source_0/N_1200 ), .C(
        \data_source_0/N_1160 ), .Y(
        \data_source_0/tag_control_sig_2_0_6[5] ));
    DFN1C0 \modulator_0/counter[4]  (.D(\modulator_0/counter_n4 ), 
        .CLK(main_clock_0_clock_out), .CLR(reset_c), .Q(
        \modulator_0/counter[4]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_16[9]  (.A(
        \data_source_0/N_1209 ), .B(\data_source_0/N_1180 ), .Y(
        \data_source_0/N_965 ));
    AO1 \data_source_0/tag_control_sig_RNO_15[6]  (.A(
        \data_source_0/N_1201 ), .B(\data_source_0/N_1173 ), .C(
        \data_source_0/N_924 ), .Y(
        \data_source_0/tag_control_sig_2_0_0[6] ));
    NOR2B \switching_circuit_0/un170_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[17] ), .B(
        main_clock_0_clock_out), .Y(
        \switching_circuit_0/un170_out_signal_switch_0_net_1 ));
    OR2 \data_source_0/counter_RNIGO4T[2]  (.A(
        \data_source_0/counter_i_0[2] ), .B(\data_source_0/N_31 ), .Y(
        \data_source_0/N_32 ));
    OR3 \data_source_0/tag_control_sig_RNO_1[7]  (.A(
        \data_source_0/tag_control_sig_2_0_0[7] ), .B(
        \data_source_0/N_936 ), .C(
        \data_source_0/tag_control_sig_2_0_8[7] ), .Y(
        \data_source_0/tag_control_sig_2_0_11[7] ));
    OR2 \data_source_0/tag_control_sig_RNO_5[16]  (.A(
        \data_source_0/N_822 ), .B(\data_source_0/N_1072 ), .Y(
        \data_source_0/tag_control_sig_2_0_2[16] ));
    AX1C \modulator_0/clock_counter_RNO[15]  (.A(AND2_0_Y), .B(
        \modulator_0/clock_counter[15]_net_1 ), .C(\modulator_0/N_89 ), 
        .Y(\modulator_0/clock_counter_n15 ));
    NOR2B \data_source_0/tag_data_buf_20_RNIAOSM[7]  (.A(
        \data_source_0/tag_data_buf_20[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[19] ));
    OR3 \data_source_0/tag_control_sig_RNO_5[11]  (.A(
        \data_source_0/N_988 ), .B(\data_source_0/N_987 ), .C(
        \data_source_0/tag_control_sig_2_0_4[11]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_12[11] ));
    OR3 \data_source_0/tag_control_sig_RNO_0[2]  (.A(
        \data_source_0/tag_control_sig_2_0_0[2] ), .B(
        \data_source_0/N_859 ), .C(
        \data_source_0/tag_control_sig_2_0_7[2] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[2] ));
    NOR2B \modulator_0/clock_counter_RNIKM0A[7]  (.A(
        \modulator_0/clock_counter_c6 ), .B(
        \modulator_0/clock_counter[7]_net_1 ), .Y(
        \modulator_0/clock_counter_c7 ));
    NOR2B \data_source_0/tag_data_buf_11_RNO[6]  (.A(
        \data_source_0/tag_data_buf_11[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_11_4[6] ));
    NOR2B \data_source_0/tag_data_buf_12_RNO[7]  (.A(
        \data_source_0/tag_data_buf_12[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_12_4[7] ));
    NOR3C \modulator_0/output_signal_RNO_0  (.A(
        \modulator_0/clock_counter[13]_net_1 ), .B(
        \modulator_0/clock_counter[15]_net_1 ), .C(
        \modulator_0/clock_counter[14]_net_1 ), .Y(
        \modulator_0/un6lto15_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_18[15]  (.A(
        \data_source_0/N_1192 ), .B(\data_source_0/N_1159 ), .Y(
        \data_source_0/N_1061 ));
    DFN1E1C0 \data_source_0/tag_data_buf_3[4]  (.D(
        \data_source_0/tag_data_buf_3_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_3[4]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_16_RNO[5]  (.A(
        \data_source_0/tag_data_buf_16[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_16_4[5] ));
    XOR2 \data_source_0/data_index_RNI3LP8[0]  (.A(
        \data_source_0/data_index[3]_net_1 ), .B(
        \data_source_0/data_index[0]_net_1 ), .Y(\data_source_0/N_748 )
        );
    NOR2B \modulator_0/counter_RNO[4]  (.A(
        \modulator_0/counter_0_sqmuxa ), .B(
        \modulator_0/counter_n4_tz ), .Y(\modulator_0/counter_n4 ));
    AND3 \data_source_0/un3_data_index_I_18  (.A(
        \data_source_0/data_index[3]_net_1 ), .B(
        \data_source_0/data_index_0[4]_net_1 ), .C(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/DWACT_FINC_E[2] ));
    NOR3B \data_source_0/tag_control_sig_RNO_14[9]  (.A(
        \data_source_0/N_1136 ), .B(
        \data_source_0/tag_control_sig_2_0_a20_3_2[9] ), .C(
        \data_source_0/N_703_i ), .Y(\data_source_0/N_960 ));
    OR3 \data_source_0/tag_control_sig_RNO[3]  (.A(
        \data_source_0/tag_control_sig_2_0_10[3] ), .B(
        \data_source_0/tag_control_sig_2_0_9[3] ), .C(
        \data_source_0/tag_control_sig_2_0_14[3] ), .Y(
        \data_source_0/tag_control_sig_2[3] ));
    OR2A \data_source_0/tag_data_buf_20_RNO[2]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_20[1]_net_1 ), .Y(
        \data_source_0/tag_data_buf_20_4[2] ));
    NOR2B \data_source_0/tag_data_buf_17_RNO[7]  (.A(
        \data_source_0/tag_data_buf_17[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_17_4[7] ));
    DFN1E1 \data_source_0/tag_control_sig[9]  (.D(
        \data_source_0/tag_control_sig_2[9] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[9] ));
    NOR2A \data_source_0/data_index_RNI7I6D[4]  (.A(
        \data_source_0/N_1133 ), .B(
        \data_source_0/data_index[4]_net_1 ), .Y(
        \data_source_0/N_1230 ));
    NOR3B \data_source_0/data_index_RNIIMJH[3]  (.A(
        \data_source_0/data_index[3]_net_1 ), .B(
        \data_source_0/tag_control_sig_1_649_3 ), .C(
        \data_source_0/data_index[6]_net_1 ), .Y(
        \data_source_0/tag_control_sig_1_649_5 ));
    NOR2B \switching_circuit_0/un30_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[3] ), .B(main_clock_0_clock_out)
        , .Y(\switching_circuit_0/un30_out_signal_switch_0_net_1 ));
    OR2A \data_source_0/tag_data_buf_4_RNO[2]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_4[1]_net_1 ), .Y(
        \data_source_0/tag_data_buf_4_4[2] ));
    NOR2B \data_source_0/data_index_RNIIF0M[5]  (.A(
        \data_source_0/N_1150 ), .B(\data_source_0/N_1133 ), .Y(
        \data_source_0/N_1187 ));
    NOR2B \data_source_0/tag_data_buf_5_RNO[3]  (.A(
        \data_source_0/tag_data_buf_5[2]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_5_4[3] ));
    XA1 \modulator_0/counter_RNO[3]  (.A(\modulator_0/counter_c2 ), .B(
        \modulator_0/counter[3]_net_1 ), .C(
        \modulator_0/counter_0_sqmuxa ), .Y(\modulator_0/counter_n3 ));
    DFN1C0 \modulator_0/counter[0]  (.D(\modulator_0/counter_n0 ), 
        .CLK(main_clock_0_clock_out), .CLR(reset_c), .Q(
        \modulator_0/counter[0]_net_1 ));
    NOR2 \data_source_0/tag_control_sig_RNO_17[18]  (.A(
        \data_source_0/data_index[2]_net_1 ), .B(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/N_1243 ));
    AO1 \data_source_0/tag_control_sig_RNO_6[3]  (.A(
        \data_source_0/N_808 ), .B(\data_source_0/N_1188 ), .C(
        \data_source_0/N_865 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[3] ));
    XA1A \data_source_0/counter_RNO[14]  (.A(\data_source_0/N_43 ), .B(
        \data_source_0/counter[14]_net_1 ), .C(
        modulator_0_output_signal), .Y(\data_source_0/counter_n14 ));
    AO1 \data_source_0/tag_control_sig_RNO_1[10]  (.A(
        \data_source_0/N_779 ), .B(\data_source_0/N_1204 ), .C(
        \data_source_0/tag_control_sig_2_0_0[10] ), .Y(
        \data_source_0/tag_control_sig_2_0_7[10] ));
    NOR2B \data_source_0/tag_control_sig_RNO_18[13]  (.A(
        \data_source_0/N_1215 ), .B(\data_source_0/N_1178 ), .Y(
        \data_source_0/N_1023 ));
    NOR2B \data_source_0/tag_data_buf_2_RNO[5]  (.A(
        \data_source_0/tag_data_buf_2[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_2_4[5] ));
    DFN1E1C0 \data_source_0/tag_data_buf_19[6]  (.D(
        \data_source_0/tag_data_buf_19_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_19[6]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_20[9]  (.A(
        \data_source_0/N_1196 ), .B(\data_source_0/N_1198 ), .Y(
        \data_source_0/N_967 ));
    XA1 \modulator_0/clock_counter_RNO[14]  (.A(
        \modulator_0/clock_counter_c13 ), .B(
        \modulator_0/clock_counter[14]_net_1 ), .C(AND2_0_Y), .Y(
        \modulator_0/clock_counter_n14 ));
    AO1 \data_source_0/tag_control_sig_RNO_12[7]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_4_1[7] ), .B(
        \data_source_0/tag_control_sig_2_0_a20_4_0[7] ), .C(
        \data_source_0/N_938 ), .Y(
        \data_source_0/tag_control_sig_2_0_4[7] ));
    NOR2B \data_source_0/tag_data_buf_20_RNO[6]  (.A(
        \data_source_0/tag_data_buf_20[5]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_20_4[6] ));
    NOR2B \data_source_0/data_index_RNID81C1_0[2]  (.A(
        \data_source_0/N_1202 ), .B(\data_source_0/N_1176 ), .Y(
        \data_source_0/N_886 ));
    OR2A \data_source_0/tag_data_buf_7_RNO[0]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_7[7]_net_1 ), .Y(
        \data_source_0/tag_data_buf_7_4[0] ));
    AO1 \data_source_0/tag_control_sig_RNO_9[9]  (.A(
        \data_source_0/N_1189 ), .B(\data_source_0/N_1176 ), .C(
        \data_source_0/N_965 ), .Y(
        \data_source_0/tag_control_sig_2_0_3[9] ));
    NOR2B \data_source_0/tag_control_sig_RNO_7[14]  (.A(
        \data_source_0/N_1187 ), .B(\data_source_0/N_1160 ), .Y(
        \data_source_0/N_1041 ));
    AO1 \data_source_0/tag_control_sig_RNO_3[0]  (.A(
        \data_source_0/N_1192 ), .B(\data_source_0/N_1162 ), .C(
        \data_source_0/N_822 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[0] ));
    NOR2B \data_source_0/data_index_RNIC90M[3]  (.A(
        \data_source_0/N_1234 ), .B(\data_source_0/N_1149 ), .Y(
        \data_source_0/N_853_2 ));
    NOR3C \data_source_0/counter_RNI43142[1]  (.A(
        \data_source_0/output_data_1_sqmuxa_i_a3_1 ), .B(
        \data_source_0/N_90 ), .C(
        \data_source_0/output_data_1_sqmuxa_i_a3_2 ), .Y(
        \data_source_0/output_data_1_sqmuxa_i_a3_4 ));
    NOR3C \data_source_0/tag_control_sig_RNO_16[7]  (.A(
        \data_source_0/data_index[2]_net_1 ), .B(
        \data_source_0/N_1140 ), .C(
        \data_source_0/tag_control_sig_2_0_a20_2_0[7] ), .Y(
        \data_source_0/N_930 ));
    DFN1C0 \data_source_0/data_index_0[4]  (.D(\data_source_0/I_12 ), 
        .CLK(modulator_0_output_signal), .CLR(reset_c), .Q(
        \data_source_0/data_index_0[4]_net_1 ));
    OR3 \data_source_0/tag_control_sig_RNO_2[10]  (.A(
        \data_source_0/tag_control_sig_2_0_6[10] ), .B(
        \data_source_0/tag_control_sig_2_0_5[10] ), .C(
        \data_source_0/tag_control_sig_2_0_9[10] ), .Y(
        \data_source_0/tag_control_sig_2_0_12[10] ));
    NOR2B \data_source_0/tag_data_buf_6_RNO[5]  (.A(
        \data_source_0/tag_data_buf_6[4]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_6_4[5] ));
    DFN1C0 \data_source_0/data_index[6]  (.D(\data_source_0/I_17 ), 
        .CLK(modulator_0_output_signal), .CLR(reset_c), .Q(
        \data_source_0/data_index[6]_net_1 ));
    AND3 \main_clock_0/un5_counter_1_I_16  (.A(
        \main_clock_0/DWACT_FINC_E[0] ), .B(
        \main_clock_0/DWACT_FINC_E[1] ), .C(
        \main_clock_0/counter[5]_net_1 ), .Y(\main_clock_0/N_3 ));
    DFN1E1C0 \data_source_0/output_data[15]  (.D(
        \data_source_0/output_data_23[15] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[15] ));
    NOR2B \data_source_0/data_index_RNIEIJH[5]  (.A(
        \data_source_0/N_1154 ), .B(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/N_1123_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_3[7]  (.A(
        \data_source_0/N_766 ), .B(\data_source_0/N_1182 ), .C(
        \data_source_0/N_931 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[7] ));
    DFN1E1C0 \data_source_0/tag_data_buf_17[7]  (.D(
        \data_source_0/tag_data_buf_17_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_17[7]_net_1 ));
    OA1 \data_source_0/tag_control_sig_RNO_3[19]  (.A(
        \data_source_0/N_1192 ), .B(\data_source_0/N_1209 ), .C(
        \data_source_0/N_1179 ), .Y(
        \data_source_0/tag_control_sig_RNO_3[19]_net_1 ));
    DFN1E1P0 \data_source_0/tag_data_buf_20[2]  (.D(
        \data_source_0/tag_data_buf_20_4[2] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_20[2]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_18[1]  (.A(
        \data_source_0/N_761 ), .B(\data_source_0/N_1196 ), .Y(
        \data_source_0/N_830 ));
    NOR2B \data_source_0/tag_data_buf_2_RNO[4]  (.A(
        \data_source_0/tag_data_buf_2[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_2_4[4] ));
    OR3 \data_source_0/tag_control_sig_RNO_8[19]  (.A(
        \data_source_0/N_1125 ), .B(\data_source_0/N_1117 ), .C(
        \data_source_0/tag_control_sig_2_0_1[19] ), .Y(
        \data_source_0/tag_control_sig_2_0_8[19] ));
    AND3 \main_clock_0/un5_counter_1_I_10  (.A(
        \main_clock_0/counter[0]_net_1 ), .B(
        \main_clock_0/counter[1]_net_1 ), .C(
        \main_clock_0/counter[2]_net_1 ), .Y(
        \main_clock_0/DWACT_FINC_E[0] ));
    NOR2A \data_source_0/data_index_RNI9RP8[7]  (.A(
        \data_source_0/data_index[7]_net_1 ), .B(
        \data_source_0/data_index[2]_net_1 ), .Y(
        \data_source_0/tag_control_sig_1_649_3 ));
    OR2A \data_source_0/tag_data_buf_13_RNO[0]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_13[7]_net_1 ), .Y(
        \data_source_0/tag_data_buf_13_4[0] ));
    AO1 \data_source_0/tag_control_sig_RNO_4[6]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_3_0[6] ), .B(
        \data_source_0/N_1233 ), .C(\data_source_0/N_919 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[6] ));
    NOR2B \data_source_0/tag_control_sig_RNO_16[4]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_7_0[4] ), .B(
        \data_source_0/N_1200 ), .Y(\data_source_0/N_889 ));
    DFN1C0 \data_source_0/counter[13]  (.D(\data_source_0/counter_n13 )
        , .CLK(main_clock_0_clock_out), .CLR(reset_c), .Q(
        \data_source_0/counter[13]_net_1 ));
    DFN1E1C0 \data_source_0/tag_data_buf_2[4]  (.D(
        \data_source_0/tag_data_buf_2_4[4] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_2[4]_net_1 ));
    DFN1E1P0 \data_source_0/tag_data_buf_17[0]  (.D(
        \data_source_0/tag_data_buf_17_4[0] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_17[0]_net_1 ));
    NOR3A \data_source_0/tag_control_sig_RNO_20[4]  (.A(
        \data_source_0/data_index[8]_net_1 ), .B(
        \data_source_0/data_index_0[7]_net_1 ), .C(
        \data_source_0/data_index[0]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_7_0[4] ));
    DFN1E1C0 \data_source_0/output_data[9]  (.D(
        \data_source_0/output_data_23[9] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[9] ));
    IOPAD_TRI \output_signal_pad[8]/U0/U0  (.D(
        \output_signal_pad[8]/U0/NET1 ), .E(
        \output_signal_pad[8]/U0/NET2 ), .PAD(output_signal[8]));
    NOR2B \data_source_0/tag_data_buf_4_RNO[1]  (.A(
        \data_source_0/tag_data_buf_4[0]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_4_4[1] ));
    DFN1E1C0 \data_source_0/output_data[17]  (.D(
        \data_source_0/output_data_23[17] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[17] ));
    NOR2B \data_source_0/tag_control_sig_RNO_3[12]  (.A(
        \data_source_0/N_1197 ), .B(\data_source_0/N_1178 ), .Y(
        \data_source_0/N_1015 ));
    AO1 \data_source_0/tag_control_sig_RNO_18[4]  (.A(
        \data_source_0/N_1200 ), .B(\data_source_0/N_1173 ), .C(
        \data_source_0/N_894 ), .Y(
        \data_source_0/tag_control_sig_2_0_7[4] ));
    NOR2B \data_source_0/tag_control_sig_RNO_15[16]  (.A(
        \data_source_0/N_1229 ), .B(\data_source_0/N_1160 ), .Y(
        \data_source_0/N_1078 ));
    AO1 \data_source_0/tag_control_sig_RNO_8[12]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_2_1[12] ), .B(
        \data_source_0/tag_control_sig_2_0_a20_2_0[12] ), .C(
        \data_source_0/N_873 ), .Y(
        \data_source_0/tag_control_sig_2_0_4[12] ));
    NOR2B \data_source_0/data_index_RNICN6D_1[9]  (.A(
        \data_source_0/data_index[9]_net_1 ), .B(
        \data_source_0/N_1142 ), .Y(\data_source_0/N_1160 ));
    OR3 \data_source_0/tag_control_sig_RNO_1[17]  (.A(
        \data_source_0/N_1091 ), .B(\data_source_0/N_1090 ), .C(
        \data_source_0/tag_control_sig_2_0_2[17] ), .Y(
        \data_source_0/tag_control_sig_2_0_9[17] ));
    DFN1E1C0 \data_source_0/tag_data_buf_2[0]  (.D(
        \data_source_0/output_data_23[1] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_2[0]_net_1 ));
    NOR2B \modulator_0/clock_counter_RNIJ6HC[9]  (.A(
        \modulator_0/clock_counter_c8 ), .B(\modulator_0/un6lto9 ), .Y(
        \modulator_0/clock_counter_c9 ));
    XOR2 \data_source_0/counter_RNO_0[5]  (.A(
        \data_source_0/counter[5]_net_1 ), .B(\data_source_0/N_34 ), 
        .Y(\data_source_0/N_53_i ));
    DFN1C0 \main_clock_0/counter[6]  (.D(\main_clock_0/I_17_0 ), .CLK(
        GLA), .CLR(reset_c), .Q(\main_clock_0/counter[6]_net_1 ));
    NOR3B \data_source_0/tag_control_sig_RNO_18[10]  (.A(
        \data_source_0/N_668 ), .B(
        \data_source_0/tag_control_sig_2_0_a20_5_0[10] ), .C(
        \data_source_0/data_index_0[4]_net_1 ), .Y(
        \data_source_0/N_979 ));
    NOR2B \data_source_0/tag_control_sig_RNO_5[6]  (.A(
        \data_source_0/N_726 ), .B(\data_source_0/N_1174 ), .Y(
        \data_source_0/N_915 ));
    IOPAD_TRI \output_signal_pad[4]/U0/U0  (.D(
        \output_signal_pad[4]/U0/NET1 ), .E(
        \output_signal_pad[4]/U0/NET2 ), .PAD(output_signal[4]));
    NOR2B \data_source_0/data_index_RNIIF0M_1[1]  (.A(
        \data_source_0/N_1151 ), .B(\data_source_0/N_1136 ), .Y(
        \data_source_0/N_1207 ));
    NOR2B \data_source_0/tag_control_sig_RNO_22[17]  (.A(
        \data_source_0/N_1217 ), .B(\data_source_0/N_1159 ), .Y(
        \data_source_0/N_1094 ));
    OR3 \data_source_0/tag_control_sig_RNO[13]  (.A(
        \data_source_0/tag_control_sig_2_0_15[13] ), .B(
        \data_source_0/tag_control_sig_2_0_14[13] ), .C(
        \data_source_0/tag_control_sig_2_0_16[13] ), .Y(
        \data_source_0/tag_control_sig_2[13] ));
    OR2A \data_source_0/tag_data_buf_5_RNO[2]  (.A(
        modulator_0_output_signal), .B(
        \data_source_0/tag_data_buf_5[1]_net_1 ), .Y(
        \data_source_0/tag_data_buf_5_4[2] ));
    NOR2B \data_source_0/tag_data_buf_18_RNO[7]  (.A(
        \data_source_0/tag_data_buf_18[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_18_4[7] ));
    OR3 \data_source_0/tag_control_sig_RNO_2[17]  (.A(
        \data_source_0/tag_control_sig_2_0_8[17] ), .B(
        \data_source_0/tag_control_sig_2_0_7[17] ), .C(
        \data_source_0/tag_control_sig_2_0_11[17] ), .Y(
        \data_source_0/tag_control_sig_2_0_14[17] ));
    XOR2 \data_source_0/un3_data_index_I_20  (.A(\data_source_0/N_4 ), 
        .B(\data_source_0/data_index[7]_net_1 ), .Y(
        \data_source_0/I_20 ));
    NOR3C \data_source_0/tag_control_sig_RNO_14[11]  (.A(
        \data_source_0/N_1180 ), .B(
        \data_source_0/tag_control_sig_1_3[649] ), .C(
        \data_source_0/N_1233 ), .Y(\data_source_0/N_987 ));
    NOR2B \data_source_0/data_index_RNID81C1[2]  (.A(
        \data_source_0/N_1215 ), .B(\data_source_0/N_1161 ), .Y(
        \data_source_0/N_879 ));
    AO1 \modulator_0/output_signal_RNO_3  (.A(\modulator_0/un6lt9 ), 
        .B(\modulator_0/un6lto9 ), .C(\modulator_0/un6lto10 ), .Y(
        \modulator_0/un6lt11 ));
    AO1 \data_source_0/tag_control_sig_RNO_23[17]  (.A(
        \data_source_0/N_1201 ), .B(\data_source_0/N_1174 ), .C(
        \data_source_0/N_1101 ), .Y(
        \data_source_0/tag_control_sig_2_0_5[17] ));
    OR2A \data_source_0/counter_RNI3DP13[10]  (.A(
        \data_source_0/counter[10]_net_1 ), .B(\data_source_0/N_39 ), 
        .Y(\data_source_0/N_40 ));
    NOR3C \data_source_0/tag_control_sig_RNO_6[13]  (.A(
        \data_source_0/N_1132 ), .B(\data_source_0/N_1229 ), .C(
        \data_source_0/N_1240 ), .Y(\data_source_0/N_1030 ));
    NOR3B \data_source_0/tag_control_sig_RNO_22[13]  (.A(
        \data_source_0/N_1185 ), .B(\data_source_0/N_1227 ), .C(
        \data_source_0/N_668 ), .Y(\data_source_0/N_1021 ));
    DFN1E1C0 \data_source_0/tag_data_buf_8[1]  (.D(
        \data_source_0/tag_data_buf_8_4[1] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_8[1]_net_1 ));
    OA1 \modulator_0/output_signal_RNO_2  (.A(\modulator_0/un5lto15_5 )
        , .B(\modulator_0/un5lto15_6 ), .C(AND2_0_Y), .Y(
        \modulator_0/output_signal_1_sqmuxa_0 ));
    NOR3C \data_source_0/tag_control_sig_RNO_10[3]  (.A(
        \data_source_0/data_index[3]_net_1 ), .B(
        \data_source_0/N_1145 ), .C(\data_source_0/N_1208 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_2_0[3] ));
    XAI1 \data_source_0/counter_RNO[6]  (.A(
        \data_source_0/counter_i_0[6] ), .B(\data_source_0/N_35 ), .C(
        modulator_0_output_signal), .Y(\data_source_0/N_16 ));
    DFN1E1 \data_source_0/tag_control_sig[8]  (.D(
        \data_source_0/tag_control_sig_2[8] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[8] ));
    MX2 \switching_circuit_0/out_signal_switch_1[17]  (.A(
        \switching_circuit_0/un170_out_signal_switch_0_net_1 ), .B(
        \switching_circuit_0/un173_out_signal_switch_0_net_1 ), .S(
        modulator_0_output_signal), .Y(\output_signal_c[17] ));
    NOR2B \data_source_0/tag_control_sig_RNO_23[13]  (.A(
        \data_source_0/N_1206 ), .B(\data_source_0/N_1181 ), .Y(
        \data_source_0/N_1034 ));
    NOR2B \data_source_0/tag_data_buf_18_RNO[2]  (.A(
        \data_source_0/tag_data_buf_18[1]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_18_4[2] ));
    NOR2B \data_source_0/tag_control_sig_RNO_15[17]  (.A(
        \data_source_0/N_1133 ), .B(
        \data_source_0/data_index[4]_net_1 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_4_1[17] ));
    NOR2B \data_source_0/data_index_RNIIF0M_1[2]  (.A(
        \data_source_0/N_1157 ), .B(\data_source_0/N_1134 ), .Y(
        \data_source_0/N_1197 ));
    DFN1E1C0 \modulator_0/clock_counter[12]  (.D(
        \modulator_0/clock_counter_n12 ), .CLK(main_clock_0_clock_out), 
        .CLR(reset_c), .E(\modulator_0/clock_countere ), .Q(
        \modulator_0/un6lto12 ));
    NOR2B \data_source_0/data_index_RNIAL6D[7]  (.A(
        \data_source_0/N_1132 ), .B(
        \data_source_0/data_index[7]_net_1 ), .Y(
        \data_source_0/N_1213 ));
    NOR2 \data_source_0/data_index_RNI9RP8_2[4]  (.A(
        \data_source_0/data_index[4]_net_1 ), .B(
        \data_source_0/data_index[5]_net_1 ), .Y(
        \data_source_0/tag_control_sig_1_3[649] ));
    NOR2B \switching_circuit_0/un40_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[4] ), .B(main_clock_0_clock_out)
        , .Y(\switching_circuit_0/un40_out_signal_switch_0_net_1 ));
    NOR2B \switching_circuit_0/un110_out_signal_switch_0  (.A(
        \data_source_0_tag_control_sig[11] ), .B(
        main_clock_0_clock_out), .Y(
        \switching_circuit_0/un110_out_signal_switch_0_net_1 ));
    NOR2A \data_source_0/tag_control_sig_RNO_20[10]  (.A(
        \data_source_0/N_1239 ), .B(\data_source_0/N_703_i ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_4_0[10] ));
    OA1 \data_source_0/tag_control_sig_RNO_17[16]  (.A(
        \data_source_0/N_1201 ), .B(\data_source_0/N_1226 ), .C(
        \data_source_0/N_1161 ), .Y(
        \data_source_0/tag_control_sig_RNO_17[16]_net_1 ));
    AO1 \data_source_0/tag_control_sig_RNO_7[3]  (.A(
        \data_source_0/N_757 ), .B(\data_source_0/N_1175 ), .C(
        \data_source_0/tag_control_sig_2_0_0[3] ), .Y(
        \data_source_0/tag_control_sig_2_0_8[3] ));
    NOR2B \data_source_0/tag_data_buf_14_RNO[4]  (.A(
        \data_source_0/tag_data_buf_14[3]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_14_4[4] ));
    NOR2B \data_source_0/tag_control_sig_RNO_3[16]  (.A(
        \data_source_0/N_1193 ), .B(\data_source_0/N_1195 ), .Y(
        \data_source_0/N_1080 ));
    NOR2B \data_source_0/output_data_RNO[2]  (.A(
        \data_source_0/tag_data_buf_3[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[2] ));
    DFN1E1 \data_source_0/tag_control_sig[4]  (.D(
        \data_source_0/tag_control_sig_2[4] ), .CLK(
        main_clock_0_clock_out), .E(
        \data_source_0/tag_control_sig_1_sqmuxa_net_1 ), .Q(
        \data_source_0_tag_control_sig[4] ));
    DFN1E1C0 \data_source_0/tag_data_buf_2[7]  (.D(
        \data_source_0/tag_data_buf_2_4[7] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_2[7]_net_1 ));
    NOR2B \data_source_0/tag_control_sig_RNO_22[7]  (.A(
        \data_source_0/N_1238 ), .B(\data_source_0/N_703_i ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_4_0[7] ));
    NOR2B \data_source_0/tag_control_sig_RNO_16[0]  (.A(
        \data_source_0/N_1207 ), .B(\data_source_0/N_1176 ), .Y(
        \data_source_0/N_827 ));
    AO1 \data_source_0/tag_control_sig_RNO_8[16]  (.A(
        \data_source_0/tag_control_sig_2_0_a20_1_0[16] ), .B(
        \data_source_0/N_1074_2 ), .C(\data_source_0/N_1028 ), .Y(
        \data_source_0/tag_control_sig_2_0_1[16] ));
    DFN1E1P0 \data_source_0/tag_data_buf_17[4]  (.D(
        \data_source_0/tag_data_buf_17_4[4] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_17[4]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_10_RNO[7]  (.A(
        \data_source_0/tag_data_buf_10[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_10_4[7] ));
    DFN1E1C0 \data_source_0/output_data[18]  (.D(
        \data_source_0/output_data_23[18] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[18] ));
    IOPAD_TRI \output_signal_pad[12]/U0/U0  (.D(
        \output_signal_pad[12]/U0/NET1 ), .E(
        \output_signal_pad[12]/U0/NET2 ), .PAD(output_signal[12]));
    AO1 \data_source_0/tag_control_sig_RNO_3[11]  (.A(
        \data_source_0/N_1207 ), .B(\data_source_0/N_1184 ), .C(
        \data_source_0/N_872 ), .Y(
        \data_source_0/tag_control_sig_2_0_2[11] ));
    NOR3B \data_source_0/tag_control_sig_RNO_6[0]  (.A(
        \data_source_0/data_index[9]_net_1 ), .B(
        \data_source_0/tag_control_sig_2_0_a20_0[0] ), .C(
        \data_source_0/data_index_0[7]_net_1 ), .Y(
        \data_source_0/N_811 ));
    AO1 \data_source_0/tag_control_sig_RNO_8[11]  (.A(
        \data_source_0/N_1242 ), .B(\data_source_0/N_1183 ), .C(
        \data_source_0/N_993 ), .Y(
        \data_source_0/tag_control_sig_2_0_9[11] ));
    XA1A \data_source_0/tag_control_sig_RNO_10[19]  (.A(
        \data_source_0/data_index[2]_net_1 ), .B(
        \data_source_0/data_index[6]_net_1 ), .C(
        \data_source_0/N_1182 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_1_0[19] ));
    NOR3C \modulator_0/counter_RNIN4AV2[4]  (.A(
        \modulator_0/counter19_0 ), .B(\modulator_0/counter19_3 ), .C(
        \modulator_0/counter19_1 ), .Y(\modulator_0/counter19 ));
    NOR2B \data_source_0/tag_control_sig_RNO_21[19]  (.A(
        \data_source_0/N_1142 ), .B(\data_source_0/N_1183 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_12_0[19] ));
    AND3 \data_source_0/un3_data_index_I_10  (.A(
        \data_source_0/data_index[0]_net_1 ), .B(
        \data_source_0/data_index[1]_net_1 ), .C(
        \data_source_0/data_index[2]_net_1 ), .Y(
        \data_source_0/DWACT_FINC_E[0] ));
    NOR3B \data_source_0/counter_RNIR35T[2]  (.A(
        \data_source_0/counter_i_0[3] ), .B(
        \data_source_0/counter_i_0[2] ), .C(
        \data_source_0/counter[9]_net_1 ), .Y(
        \data_source_0/output_data_1_sqmuxa_i_a3_2 ));
    IOTRI_OB_EB \output_signal_pad[17]/U0/U1  (.D(
        \output_signal_c[17] ), .E(VCC), .DOUT(
        \output_signal_pad[17]/U0/NET1 ), .EOUT(
        \output_signal_pad[17]/U0/NET2 ));
    DFN1E1C0 \data_source_0/tag_data_buf_10[6]  (.D(
        \data_source_0/tag_data_buf_10_4[6] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_10[6]_net_1 ));
    NOR2A \data_source_0/tag_control_sig_RNO_24[18]  (.A(
        \data_source_0/N_1176 ), .B(\data_source_0/N_701_i ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_4_0[18] ));
    IOIN_IB \mac_control_signal_pad/U0/U1  (.YIN(
        \mac_control_signal_pad/U0/NET1 ), .Y(mac_control_signal_c));
    OR3 \data_source_0/tag_control_sig_RNO_1[18]  (.A(
        \data_source_0/N_1110 ), .B(\data_source_0/N_886 ), .C(
        \data_source_0/tag_control_sig_2_0_2[18] ), .Y(
        \data_source_0/tag_control_sig_2_0_9[18] ));
    DFN1E1C0 \data_source_0/tag_data_buf_4[1]  (.D(
        \data_source_0/tag_data_buf_4_4[1] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_4[1]_net_1 ));
    NOR2B \data_source_0/tag_data_buf_10_RNI9KMI[7]  (.A(
        \data_source_0/tag_data_buf_10[7]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/output_data_23[9] ));
    DFN1E1P0 \data_source_0/tag_data_buf_19[0]  (.D(
        \data_source_0/tag_data_buf_19_4[0] ), .CLK(
        main_clock_0_clock_out), .PRE(reset_c), .E(
        \data_source_0/N_29 ), .Q(
        \data_source_0/tag_data_buf_19[0]_net_1 ));
    XA1A \switching_circuit_0/un143_out_signal_switch_0  (.A(
        main_clock_0_clock_out), .B(\data_source_0_output_data_0[14] ), 
        .C(\data_source_0_tag_control_sig[14] ), .Y(
        \switching_circuit_0/un143_out_signal_switch_0_net_1 ));
    NOR2B \data_source_0/tag_data_buf_6_RNO[7]  (.A(
        \data_source_0/tag_data_buf_6[6]_net_1 ), .B(
        modulator_0_output_signal), .Y(
        \data_source_0/tag_data_buf_6_4[7] ));
    NOR2B \data_source_0/tag_control_sig_RNO_21[16]  (.A(
        \data_source_0/N_1152 ), .B(\data_source_0/N_1159 ), .Y(
        \data_source_0/tag_control_sig_2_0_a20_4_0[16] ));
    DFN1E1C0 \data_source_0/output_data[5]  (.D(
        \data_source_0/output_data_23[5] ), .CLK(
        main_clock_0_clock_out), .CLR(reset_c), .E(
        \data_source_0/N_29 ), .Q(\data_source_0_output_data_0[5] ));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
